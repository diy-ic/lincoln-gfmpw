* NGSPICE file created from ram_6x64.ext - technology: gf180mcuD

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_2 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_4 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_12 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_8 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_4 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_4 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_4 I0 I1 I2 I3 S0 S1 Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_2 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_4 I ZN VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VNW VPW VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_12 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_12 I Z VDD VNW VPW VSS
.ends

.subckt ram_6x64 address_i[0] address_i[1] address_i[2] address_i[3] address_i[4]
+ address_i[5] clk_i data_i[0] data_i[10] data_i[11] data_i[12] data_i[13] data_i[14]
+ data_i[15] data_i[16] data_i[17] data_i[18] data_i[19] data_i[1] data_i[20] data_i[21]
+ data_i[22] data_i[23] data_i[24] data_i[25] data_i[26] data_i[27] data_i[28] data_i[29]
+ data_i[2] data_i[30] data_i[31] data_i[3] data_i[4] data_i[5] data_i[6] data_i[7]
+ data_i[8] data_i[9] data_o[0] data_o[10] data_o[11] data_o[12] data_o[13] data_o[14]
+ data_o[15] data_o[16] data_o[17] data_o[18] data_o[19] data_o[1] data_o[20] data_o[21]
+ data_o[22] data_o[23] data_o[24] data_o[25] data_o[26] data_o[27] data_o[28] data_o[29]
+ data_o[2] data_o[30] data_o[31] data_o[3] data_o[4] data_o[5] data_o[6] data_o[7]
+ data_o[8] data_o[9] vdd vss we_i
X_06883_ _03113_ _03114_ _03115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
X_09671_ _04699_ _01998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08622_ _04114_ _01534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_85_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08553_ _04077_ _01502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08334__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07504_ memory\[59\]\[9\] _03327_ _03493_ _03503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11094__A1 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08484_ _03758_ memory\[21\]\[3\] _04037_ _04041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10141__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_175_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07435_ _03465_ _00996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10249__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12665__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07366_ _03427_ _00965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09105_ _04233_ memory\[2\]\[24\] _04380_ _04385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07297_ memory\[11\]\[10\] _03329_ _03390_ _03391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13218__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09036_ _04348_ _01714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09974__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10913__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12441__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07494__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13509__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11808__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09938_ _04842_ _00042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_142_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_142_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09869_ _04606_ memory\[40\]\[15\] _04800_ _04806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08573__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11900_ memory\[46\]\[5\] memory\[47\]\[5\] _05907_ _06111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12880_ memory\[46\]\[19\] memory\[47\]\[19\] _06596_ _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09214__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11831_ _05741_ _06042_ _06043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12639__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11543__I _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14550_ _01589_ clknet_leaf_82_clk_i memory\[24\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11762_ memory\[46\]\[3\] memory\[47\]\[3\] _05907_ _05975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13501_ memory\[62\]\[29\] memory\[63\]\[29\] _02448_ _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10713_ _05268_ _00391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14481_ _01520_ clknet_leaf_103_clk_i memory\[22\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10683__I1 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11693_ _05701_ _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_138_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13432_ _02358_ _02815_ _02822_ _02823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_192_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10644_ memory\[51\]\[12\] _03162_ _05229_ _05232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12585__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13363_ _02754_ _02755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10575_ _05031_ memory\[50\]\[12\] _05192_ _05195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_118_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15102_ _00061_ clknet_leaf_440_clk_i memory\[42\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09884__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12314_ memory\[8\]\[11\] memory\[9\]\[11\] memory\[10\]\[11\] memory\[11\]\[11\]
+ _05893_ _06032_ _06519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_134_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13294_ memory\[30\]\[25\] memory\[31\]\[25\] _02084_ _02687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15033_ _02072_ clknet_leaf_55_clk_i memory\[3\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10823__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12245_ memory\[38\]\[10\] memory\[39\]\[10\] _06039_ _06451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_114_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10199__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12176_ memory\[32\]\[9\] memory\[33\]\[9\] memory\[34\]\[9\] memory\[35\]\[9\] _06314_
+ _05743_ _06383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_120_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11127_ _03340_ memory\[58\]\[15\] _05482_ _05488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11058_ _05451_ _00553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08564__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10009_ _04610_ memory\[42\]\[17\] _04872_ _04880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10371__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14817_ _01856_ clknet_leaf_426_clk_i memory\[33\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13154__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12549__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15797_ _00756_ clknet_leaf_58_clk_i net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08316__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14748_ _01787_ clknet_leaf_391_clk_i memory\[31\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08963__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12485__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14679_ _01718_ clknet_leaf_85_clk_i memory\[28\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_79 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09858__I _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07220_ memory\[39\]\[15\] _03340_ _03330_ _03341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_15_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08619__I1 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_133_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07151_ _03200_ memory\[13\]\[24\] _03290_ _03295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07082_ _03203_ memory\[16\]\[25\] _03251_ _03257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12328__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10733__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07055__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07984_ _03762_ memory\[12\]\[5\] _03752_ _03763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08002__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09723_ _04727_ _02022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06935_ _03125_ _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12500__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_58_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09654_ _04598_ memory\[37\]\[11\] _04689_ _04691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10362__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08605_ _04104_ _01527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09585_ _04654_ _01957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08307__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08536_ _03810_ memory\[21\]\[28\] _04059_ _04068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10114__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__I1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08467_ _04031_ _01462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10908__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07530__I1 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07418_ memory\[49\]\[1\] _03311_ _03455_ _03457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08398_ _03808_ memory\[1\]\[27\] _03987_ _03995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07349_ _03418_ _00957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_5_6__f_clk_i clknet_2_0_0_clk_i clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_98_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10707__I _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10360_ _05020_ memory\[47\]\[7\] _05073_ _05081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_115_Left_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_115_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09019_ _04339_ _01706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10291_ _05036_ _00201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_76_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13611__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07046__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12030_ _05699_ _06231_ _06238_ _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09209__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13239__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_335_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11538__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07952__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13981_ _01020_ clknet_leaf_333_clk_i memory\[59\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08546__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15720_ _00679_ clknet_leaf_237_clk_i memory\[61\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12932_ memory\[14\]\[20\] memory\[15\]\[20\] _02193_ _02330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_124_Left_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15651_ _00610_ clknet_leaf_312_clk_i memory\[5\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12863_ memory\[12\]\[19\] memory\[13\]\[19\] _06714_ _02262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13047__A2 _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11273__I _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14602_ _01641_ clknet_leaf_186_clk_i memory\[26\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11814_ memory\[12\]\[4\] memory\[13\]\[4\] _06025_ _06026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08783__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15582_ _00541_ clknet_leaf_326_clk_i memory\[57\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12794_ memory\[14\]\[18\] memory\[15\]\[18\] _02193_ _02194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14533_ _01572_ clknet_leaf_360_clk_i memory\[24\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11745_ memory\[12\]\[3\] memory\[13\]\[3\] _05716_ _05958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10656__I1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07521__I1 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_155_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_155_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14464_ _01503_ clknet_leaf_352_clk_i memory\[22\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11676_ _05889_ _05890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_154_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13415_ _02216_ _02805_ _02806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10627_ memory\[51\]\[4\] _03137_ _05218_ _05223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_172_3694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14395_ _01434_ clknet_leaf_395_clk_i memory\[1\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_133_Left_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_3_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11230__A1 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13346_ _02337_ _02733_ _02735_ _02737_ _02738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10558_ _05014_ memory\[50\]\[4\] _05181_ _05186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13277_ memory\[36\]\[25\] memory\[37\]\[25\] _02338_ _02670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10489_ _05149_ _00286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15016_ _02055_ clknet_leaf_250_clk_i memory\[3\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09119__S _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12228_ memory\[0\]\[10\] memory\[1\]\[10\] memory\[2\]\[10\] memory\[3\]\[10\] _06020_
+ _06090_ _06434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11448__I _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12159_ memory\[6\]\[9\] memory\[7\]\[9\] _05706_ _06366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08958__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10592__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_142_Left_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08757__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12279__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_56_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09789__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08693__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09370_ _04525_ _01871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08321_ _03954_ _01393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08252_ _03798_ memory\[17\]\[22\] _03915_ _03918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_151_Left_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_284_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07203_ _03155_ _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08183_ _03881_ _01328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07134_ _03175_ memory\[13\]\[16\] _03279_ _03286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_6_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07065_ _03178_ memory\[16\]\[17\] _03240_ _03248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09029__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12721__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08776__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10583__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_160_Left_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_96_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input36_I data_i[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07772__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07967_ _03115_ _03750_ _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_96_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08528__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11294__S _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09706_ _04718_ _02014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06918_ _03143_ _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07898_ _03129_ memory\[19\]\[1\] _03711_ _03713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09637_ _04581_ memory\[37\]\[3\] _04678_ _04682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_28__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09699__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09568_ _04645_ _01949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08519_ _04036_ _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_33_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09499_ _04599_ _01926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11530_ _05732_ _05735_ _05740_ _05745_ _05746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_92_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_137_Right_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11461_ _03120_ _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XTAP_TAPCELL_ROW_78_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13200_ _02593_ _02594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10412_ _03227_ _03451_ _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_11392_ _03332_ memory\[62\]\[11\] _05627_ _05629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14180_ _01219_ clknet_leaf_338_clk_i memory\[19\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11469__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13131_ _06835_ _02525_ _02178_ _02526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10343_ _05071_ _00218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10373__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_131_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10274_ _05024_ memory\[46\]\[9\] _05006_ _05025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13062_ memory\[48\]\[22\] memory\[49\]\[22\] memory\[50\]\[22\] memory\[51\]\[22\]
+ _06699_ _06839_ _02458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_103_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08767__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12712__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12013_ _06149_ _06221_ _06222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07682__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_191_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13964_ _01003_ clknet_leaf_258_clk_i memory\[49\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_109_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15703_ _00662_ clknet_leaf_149_clk_i memory\[60\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12915_ memory\[54\]\[20\] memory\[55\]\[20\] _02312_ _02313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13895_ _00934_ clknet_leaf_212_clk_i memory\[11\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15634_ _00593_ clknet_leaf_163_clk_i memory\[58\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_17_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12846_ _02170_ _02244_ _02245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_158_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_17_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12779__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15565_ _00524_ clknet_leaf_228_clk_i memory\[56\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10629__I1 _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12777_ memory\[54\]\[18\] memory\[55\]\[18\] _06421_ _02177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14516_ _01555_ clknet_leaf_105_clk_i memory\[23\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11728_ _05668_ _05940_ _05941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08018__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15496_ _00455_ clknet_leaf_290_clk_i memory\[54\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14447_ _01486_ clknet_leaf_188_clk_i memory\[21\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_104_Right_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_154_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11659_ _05654_ _05867_ _05870_ _05872_ _05873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_181_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07857__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14378_ _01417_ clknet_leaf_170_clk_i memory\[1\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11379__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13329_ memory\[0\]\[26\] memory\[1\]\[26\] memory\[2\]\[26\] memory\[3\]\[26\] _05784_
+ _03226_ _02721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_0_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12703__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08758__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13594__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08870_ _04260_ _01636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07592__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07821_ _03671_ _01176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_402_clk_i clknet_5_3__leaf_clk_i clknet_leaf_402_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07752_ _03215_ memory\[63\]\[29\] _03625_ _03635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12003__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09183__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07683_ _03598_ _01111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12482__A3 _06669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_56_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09422_ _04210_ memory\[34\]\[13\] _04549_ _04553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11690__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06936__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_417_clk_i clknet_5_2__leaf_clk_i clknet_leaf_417_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12314__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09353_ _04516_ _01863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08304_ _03945_ _01385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10245__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09284_ _04208_ memory\[32\]\[12\] _04477_ _04480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_24__f_clk_i clknet_2_3_0_clk_i clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08235_ _03781_ memory\[17\]\[14\] _03904_ _03909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12673__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08166_ _03872_ _01320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11797__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08997__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07117_ _03150_ memory\[13\]\[8\] _03268_ _03277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08097_ _03781_ memory\[15\]\[14\] _03830_ _03835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09982__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07048_ _03153_ memory\[16\]\[9\] _03229_ _03239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13742__I0 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10921__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08598__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10556__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13517__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08999_ _04195_ memory\[28\]\[6\] _04322_ _04329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11816__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13009__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_173_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10961_ _05400_ _00507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12848__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12700_ memory\[60\]\[17\] memory\[61\]\[17\] _06273_ _02101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13680_ _05753_ _03066_ _05687_ _03067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11681__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10892_ memory\[55\]\[0\] _03110_ _05363_ _05364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09222__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12631_ _05675_ _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_191_4045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_4056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11551__I _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15350_ _00309_ clknet_leaf_150_clk_i memory\[4\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12562_ _06276_ _06762_ _06690_ _06763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_152_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14301_ _01340_ clknet_leaf_366_clk_i memory\[17\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13679__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11513_ _05715_ _05718_ _05723_ _05728_ _05729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15281_ _00240_ clknet_leaf_43_clk_i memory\[47\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12493_ memory\[52\]\[14\] memory\[53\]\[14\] _06143_ _06695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14232_ _01271_ clknet_leaf_138_clk_i memory\[12\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11444_ _05659_ _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_150_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12933__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11199__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13281__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14163_ _01202_ clknet_leaf_119_clk_i memory\[7\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11375_ _03315_ memory\[62\]\[3\] _05616_ _05620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09892__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13114_ memory\[16\]\[22\] memory\[17\]\[22\] memory\[18\]\[22\] memory\[19\]\[22\]
+ _02233_ _02376_ _02510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_104_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10326_ _03205_ _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_14094_ _01133_ clknet_leaf_219_clk_i memory\[63\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13045_ _02367_ _02437_ _02439_ _02441_ _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_167_3582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10831__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10257_ _05013_ _00190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_167_3593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_232_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08301__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10188_ _04585_ memory\[45\]\[5\] _04969_ _04975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_128_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14996_ _02035_ clknet_leaf_66_clk_i memory\[38\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09165__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12544__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13947_ _00986_ clknet_leaf_387_clk_i memory\[8\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11662__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xload_slew74 net75 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_159_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13878_ _00917_ clknet_leaf_66_clk_i memory\[39\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15617_ _00576_ clknet_leaf_324_clk_i memory\[58\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12829_ memory\[20\]\[18\] memory\[21\]\[18\] _06477_ _02229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10278__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11461__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15548_ _00507_ clknet_leaf_328_clk_i memory\[56\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08971__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15479_ _00438_ clknet_leaf_267_clk_i memory\[53\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12493__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08020_ _03177_ _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_141_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12506__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08979__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10786__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07651__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09971_ _04859_ _00058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12527__I1 memory\[39\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08922_ _04288_ _01660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10741__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10538__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_341_clk_i clknet_5_9__leaf_clk_i clknet_leaf_341_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09307__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08853_ _04185_ memory\[26\]\[1\] _04250_ _04252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07804_ _03191_ memory\[6\]\[21\] _03661_ _03663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08784_ _04205_ _01605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09156__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07735_ _03626_ _01135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08903__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_356_clk_i clknet_5_8__leaf_clk_i clknet_leaf_356_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11663__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07666_ _03187_ memory\[10\]\[20\] _03589_ _03590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_434_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10710__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09405_ _04193_ memory\[34\]\[5\] _04538_ _04544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10188__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07597_ _03187_ memory\[0\]\[20\] _03552_ _03553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09336_ _04507_ _01855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13499__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09267_ _04191_ memory\[32\]\[4\] _04466_ _04471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_181_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08218_ _03764_ memory\[17\]\[6\] _03893_ _03900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07890__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09198_ _04434_ _01790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08149_ _03863_ _01312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07296__I _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11160_ _03373_ memory\[58\]\[31\] _05470_ _05505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07642__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11747__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13715__I0 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10111_ _04934_ _00123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11091_ _05468_ _00569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_8_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_309_clk_i clknet_5_14__leaf_clk_i clknet_leaf_309_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09395__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10042_ _04573_ memory\[43\]\[0\] _04897_ _04898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_output67_I net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11546__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14850_ _01889_ clknet_leaf_430_clk_i memory\[34\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07960__S _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13801_ _00840_ clknet_leaf_208_clk_i memory\[16\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_162_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14781_ _01820_ clknet_leaf_428_clk_i memory\[32\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11993_ _05788_ _06202_ _05792_ _06203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_193_4107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13732_ _03350_ memory\[9\]\[20\] _03097_ _03098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10944_ memory\[55\]\[25\] _03202_ _05385_ _05391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10701__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13663_ _03049_ _03050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10098__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10875_ _05058_ memory\[54\]\[25\] _05348_ _05354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15402_ _00361_ clknet_leaf_238_clk_i memory\[51\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12614_ memory\[22\]\[15\] memory\[23\]\[15\] _06751_ _06815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13594_ memory\[38\]\[30\] memory\[39\]\[30\] _05662_ _02982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15333_ _00292_ clknet_leaf_312_clk_i memory\[4\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12545_ _06610_ _06746_ _06747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15264_ _00223_ clknet_leaf_417_clk_i memory\[47\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12476_ memory\[22\]\[13\] memory\[23\]\[13\] _06062_ _06679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14215_ _01254_ clknet_leaf_202_clk_i memory\[12\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11427_ _03367_ memory\[62\]\[28\] _05638_ _05647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_169_3622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15195_ _00154_ clknet_leaf_0_clk_i memory\[44\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14146_ _01185_ clknet_leaf_300_clk_i memory\[7\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11358_ _05610_ _00694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13006__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13706__I0 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10309_ _05047_ memory\[46\]\[20\] _05048_ _05049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14077_ _01116_ clknet_leaf_311_clk_i memory\[63\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11289_ _05573_ _00662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_383_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13331__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09127__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13182__I1 net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13028_ memory\[40\]\[21\] memory\[41\]\[21\] memory\[42\]\[21\] memory\[43\]\[21\]
+ _06875_ _02217_ _02425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08031__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11193__I0 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07870__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11392__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14979_ _02018_ clknet_leaf_403_clk_i memory\[38\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07520_ _03511_ _01035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07451_ memory\[49\]\[17\] _03344_ _03466_ _03474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13398__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09797__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07382_ _03435_ _00973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_88_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09121_ _03124_ _03855_ _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_161_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12070__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13112__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09052_ _04356_ _01722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07872__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08206__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08003_ _03775_ memory\[12\]\[11\] _03773_ _03776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12951__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10759__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_637 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1088 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07624__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08005__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_280_clk_i clknet_5_12__leaf_clk_i clknet_leaf_280_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09954_ _04623_ memory\[41\]\[23\] _04847_ _04851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09037__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13322__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09377__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12756__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08905_ _04237_ memory\[26\]\[26\] _04272_ _04279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_5_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09885_ _04814_ _00017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10270__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_128_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08836_ _04240_ _01622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08876__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09129__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12508__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07552__A2 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_295_clk_i clknet_5_15__leaf_clk_i clknet_leaf_295_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08767_ _04193_ memory\[25\]\[5\] _04183_ _04194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07718_ _03617_ _01127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08698_ _04154_ _01570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_64_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07649_ _03163_ memory\[10\]\[12\] _03578_ _03581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_64_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10660_ _05217_ _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_81_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09301__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09319_ _04243_ memory\[32\]\[29\] _04488_ _04498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10646__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10591_ _05180_ _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_69_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12330_ _06325_ _06534_ _06535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_233_clk_i clknet_5_15__leaf_clk_i clknet_leaf_233_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07863__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12261_ _03224_ _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_121_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14000_ _01039_ clknet_leaf_177_clk_i memory\[59\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_146_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11212_ _03357_ memory\[5\]\[23\] _05529_ _05533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07615__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12192_ _05921_ _06398_ _06399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_102_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput42 net42 data_o[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_147_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_248_clk_i clknet_5_27__leaf_clk_i clknet_leaf_248_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xoutput53 net53 data_o[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11143_ _05496_ _00593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10381__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput64 net64 data_o[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_164_3530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13313__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11074_ _05052_ memory\[57\]\[22\] _05457_ _05460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13692__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08040__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10025_ _04888_ _00083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14902_ _01941_ clknet_leaf_72_clk_i memory\[35\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08786__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14833_ _01872_ clknet_leaf_61_clk_i memory\[33\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12419__A3 _06602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14764_ _01803_ clknet_leaf_126_clk_i memory\[31\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11976_ _05691_ _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_114_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13715_ _03334_ memory\[9\]\[12\] _03086_ _03089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10927_ memory\[55\]\[17\] _03177_ _05374_ _05382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14695_ _01734_ clknet_5_25__leaf_clk_i memory\[2\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13646_ _05747_ _03028_ _03030_ _03032_ _03033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_128_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10858_ _05041_ memory\[54\]\[17\] _05337_ _05345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12052__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10556__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13577_ memory\[4\]\[30\] memory\[5\]\[30\] _05789_ _02965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10789_ _05308_ _00427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10989__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15316_ _00275_ clknet_leaf_263_clk_i memory\[48\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12528_ _06450_ _06729_ _06177_ _06730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11650__I1 net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12056__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15247_ _00206_ clknet_leaf_273_clk_i memory\[46\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12459_ memory\[44\]\[13\] memory\[45\]\[13\] _06319_ _06662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07865__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_1_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15178_ _00137_ clknet_leaf_38_clk_i memory\[44\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_184_3917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11387__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14129_ _01168_ clknet_leaf_123_clk_i memory\[6\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11953__I2 memory\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13304__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06951_ _03168_ _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11166__I0 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08031__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12902__I1 net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11866__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09670_ _04614_ memory\[37\]\[19\] _04689_ _04699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06882_ net5 net6 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XFILLER_0_94_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_19_Left_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_27_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08621_ memory\[23\]\[3\] _03315_ _04110_ _04114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_85_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08552_ _03758_ memory\[22\]\[3\] _04073_ _04077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11618__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07105__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07503_ _03502_ _01027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08483_ _04040_ _01469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12291__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07434_ memory\[49\]\[9\] _03327_ _03455_ _03465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06944__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12043__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13350__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07365_ _03156_ memory\[8\]\[10\] _03426_ _03427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10466__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_28_Left_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_165_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09104_ _04384_ _01746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07296_ _03378_ _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_5_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_54_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13218__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09035_ _04231_ memory\[28\]\[23\] _04344_ _04348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09598__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13543__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08270__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09990__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09937_ _04606_ memory\[41\]\[15\] _04836_ _04842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_37_Left_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_42_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_279_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_142_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09868_ _04805_ _00009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08819_ _03193_ _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09799_ memory\[3\]\[15\] _03171_ _04762_ _04768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13017__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11830_ memory\[32\]\[4\] memory\[33\]\[4\] memory\[34\]\[4\] memory\[35\]\[4\] _05742_
+ _05743_ _06042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11609__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06918__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09522__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11761_ _05973_ _05974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12856__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11760__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_331_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13500_ _02888_ _02889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10712_ _05031_ memory\[52\]\[12\] _05265_ _05268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14480_ _01519_ clknet_leaf_101_clk_i memory\[22\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11692_ _05905_ _05906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_181_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Left_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09230__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13431_ _02367_ _02817_ _02819_ _02821_ _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08089__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_172_clk_i clknet_5_28__leaf_clk_i clknet_leaf_172_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12034__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10643_ _05231_ _00358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13362_ memory\[20\]\[26\] memory\[21\]\[26\] _02368_ _02754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07836__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10574_ _05194_ _00326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_118_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15101_ _00060_ clknet_leaf_434_clk_i memory\[42\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12313_ _06028_ _06517_ _06304_ _06518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_13293_ _02685_ _02686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_121_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_187_clk_i clknet_5_29__leaf_clk_i clknet_leaf_187_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_146_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15032_ _02071_ clknet_leaf_59_clk_i memory\[3\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12244_ _05659_ _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11396__I0 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12175_ _05736_ _06381_ _06177_ _06382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_20_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11126_ _05487_ _00585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_110_clk_i clknet_5_22__leaf_clk_i clknet_leaf_110_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11148__I0 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11057_ _05035_ memory\[57\]\[14\] _05446_ _05451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09405__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09761__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10008_ _04879_ _00075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_125_clk_i clknet_5_29__leaf_clk_i clknet_leaf_125_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14816_ _01855_ clknet_leaf_420_clk_i memory\[33\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15796_ _00755_ clknet_leaf_58_clk_i net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13065__A3 _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09513__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14747_ _01786_ clknet_leaf_0_clk_i memory\[30\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11959_ _06028_ _06168_ _05722_ _06169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_87_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11670__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14678_ _01717_ clknet_leaf_84_clk_i memory\[28\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_104_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13629_ memory\[56\]\[31\] memory\[57\]\[31\] memory\[58\]\[31\] memory\[59\]\[31\]
+ _05711_ _03748_ _03016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_15_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__I1 _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07150_ _03294_ _00882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07081_ _03256_ _00851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12328__A2 _06532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11387__I0 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_39_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08252__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07983_ _03140_ _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_96_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_280_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09722_ _04598_ memory\[38\]\[11\] _04725_ _04727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06934_ _03155_ _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11839__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13384__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09315__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09653_ _04690_ _01989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_18__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08604_ _03810_ memory\[22\]\[28\] _04095_ _04104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09584_ _04595_ memory\[36\]\[10\] _04653_ _04654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_26_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09504__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_118_Right_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08535_ _04067_ _01494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08466_ _03808_ memory\[20\]\[27\] _04023_ _04031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07417_ _03456_ _00987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10196__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08397_ _03994_ _01429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09807__I1 _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07348_ _03132_ memory\[8\]\[2\] _03415_ _03418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_98_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07294__I1 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07279_ _03381_ _00924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_59_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09018_ _04214_ memory\[28\]\[15\] _04333_ _04339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10290_ _05035_ memory\[46\]\[14\] _05027_ _05036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11819__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13611__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08243__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13119__I1 net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10050__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11755__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13980_ _01019_ clknet_leaf_328_clk_i memory\[59\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_42_clk_i clknet_5_18__leaf_clk_i clknet_leaf_42_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09743__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12931_ _02328_ _02329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12862_ _06844_ _02256_ _02258_ _02260_ _02261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15650_ _00609_ clknet_leaf_282_clk_i memory\[5\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13047__A3 _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14601_ _01640_ clknet_leaf_180_clk_i memory\[26\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11813_ _05677_ _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15581_ _00540_ clknet_leaf_333_clk_i memory\[57\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_159_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12793_ _05683_ _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_57_clk_i clknet_5_20__leaf_clk_i clknet_leaf_57_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_115_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14532_ _01571_ clknet_leaf_361_clk_i memory\[24\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11744_ _05700_ _05952_ _05954_ _05956_ _05957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_55_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12007__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14463_ _01502_ clknet_leaf_348_clk_i memory\[22\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11675_ memory\[12\]\[2\] memory\[13\]\[2\] _05716_ _05889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13414_ memory\[40\]\[27\] memory\[41\]\[27\] memory\[42\]\[27\] memory\[43\]\[27\]
+ _05692_ _02217_ _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_92_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10626_ _05222_ _00350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_172_3684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14394_ _01433_ clknet_leaf_30_clk_i memory\[1\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_172_3695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13345_ _02344_ _02736_ _02737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_10_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10557_ _05185_ _00318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11230__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13276_ _02319_ _02661_ _02668_ _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_10488_ _05012_ memory\[4\]\[3\] _05145_ _05149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11369__I0 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15015_ _02054_ clknet_leaf_251_clk_i memory\[3\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12227_ _06159_ _06432_ _06018_ _06433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_110_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09982__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12158_ _06364_ _06365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__13366__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11109_ _05478_ _00577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12089_ memory\[0\]\[8\] memory\[1\]\[8\] memory\[2\]\[8\] memory\[3\]\[8\] _06020_
+ _06090_ _06297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_34_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09135__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09734__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_91_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_152_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12246__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15779_ _00738_ clknet_leaf_336_clk_i net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08320_ _03798_ memory\[18\]\[22\] _03951_ _03954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08251_ _03917_ _01360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_227_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07202_ _03328_ _00900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08182_ _03796_ memory\[29\]\[21\] _03879_ _03881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07133_ _03285_ _00874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07276__I1 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07064_ _03247_ _00843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_12_Right_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08214__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10032__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_103_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_71_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07966_ _03749_ _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__09045__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09705_ _04581_ memory\[38\]\[3\] _04714_ _04718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input29_I data_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06917_ net35 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_74_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07897_ _03712_ _01211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09636_ _04681_ _01981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08884__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_21_Right_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12237__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09567_ _04579_ memory\[36\]\[2\] _04642_ _04645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10919__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08518_ _04058_ _01486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_137_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09498_ _04598_ memory\[35\]\[11\] _04596_ _04599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_137_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08449_ _03791_ memory\[20\]\[19\] _04012_ _04022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_34_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_108_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11460_ _05675_ _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_135_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10411_ _05107_ _00250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08464__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11391_ _05628_ _00709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10654__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_30_Right_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_150_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10271__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07967__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13130_ memory\[54\]\[23\] memory\[55\]\[23\] _02312_ _02525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10342_ _05070_ memory\[46\]\[31\] _05005_ _05071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08124__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_429_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08216__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13596__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13061_ _06835_ _02456_ _02178_ _02457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10273_ _03152_ _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_103_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12012_ memory\[48\]\[7\] memory\[49\]\[7\] memory\[50\]\[7\] memory\[51\]\[7\] _06010_
+ _06150_ _06221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11993__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09964__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_176_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13963_ _01002_ clknet_leaf_239_clk_i memory\[49\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15702_ _00661_ clknet_leaf_149_clk_i memory\[60\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12914_ _05683_ _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13894_ _00933_ clknet_leaf_216_clk_i memory\[11\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15633_ _00592_ clknet_leaf_176_clk_i memory\[58\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12845_ memory\[56\]\[19\] memory\[57\]\[19\] memory\[58\]\[19\] memory\[59\]\[19\]
+ _06827_ _02171_ _02244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_185_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_17_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10829__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15564_ _00523_ clknet_leaf_227_clk_i memory\[56\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12776_ _02175_ _02176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_115_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14515_ _01554_ clknet_leaf_100_clk_i memory\[23\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11727_ memory\[56\]\[3\] memory\[57\]\[3\] memory\[58\]\[3\] memory\[59\]\[3\] _05670_
+ _05671_ _05940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_56_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15495_ _00454_ clknet_5_15__leaf_clk_i memory\[54\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14446_ _01485_ clknet_leaf_190_clk_i memory\[21\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11658_ _05668_ _05871_ _05872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_141_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10609_ _05212_ _00343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14377_ _01416_ clknet_leaf_249_clk_i memory\[1\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10564__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11589_ memory\[60\]\[1\] memory\[61\]\[1\] _05656_ _05804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07937__I _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10262__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13328_ _05752_ _02719_ _05791_ _02720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_12_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08034__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13259_ _06838_ _02651_ _02652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08969__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07820_ _03215_ memory\[6\]\[29\] _03661_ _03671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_32_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07430__I1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09707__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07751_ _03634_ _01143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07682_ _03212_ memory\[10\]\[28\] _03589_ _03598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09421_ _04552_ _01895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12482__A4 _06684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12219__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10739__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12314__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09352_ _04208_ memory\[33\]\[12\] _04513_ _04516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08303_ _03781_ memory\[18\]\[14\] _03940_ _03945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07113__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_378_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09283_ _04479_ _01830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08234_ _03908_ _01352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06952__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08008__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08165_ _03779_ memory\[29\]\[13\] _03868_ _03872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10474__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10253__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07116_ _03276_ _00866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08096_ _03834_ _01288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_430_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10273__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07047_ _03238_ _00835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_73_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07783__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10005__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08998_ _04328_ _01696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07949_ _03739_ _01236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_170_Right_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10960_ _05004_ memory\[56\]\[0\] _05399_ _05400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09619_ _04631_ memory\[36\]\[27\] _04664_ _04672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10891_ _05362_ _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11681__A2 _05894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12630_ _06272_ _06824_ _06826_ _06829_ _06830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06926__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12561_ memory\[62\]\[15\] memory\[63\]\[15\] _06557_ _06762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07488__I1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08685__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12630__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14300_ _01339_ clknet_leaf_367_clk_i memory\[17\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07958__S _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11512_ _05724_ _05727_ _05728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_80_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15280_ _00239_ clknet_leaf_44_clk_i memory\[47\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12492_ _06272_ _06688_ _06691_ _06693_ _06694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_0_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_81_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14231_ _01270_ clknet_leaf_112_clk_i memory\[12\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08437__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11443_ _03118_ _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_34_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14162_ _01201_ clknet_leaf_119_clk_i memory\[7\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11374_ _05619_ _00701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13113_ _02371_ _02508_ _02373_ _02509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10325_ _05059_ _00212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14093_ _01132_ clknet_leaf_224_clk_i memory\[63\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13044_ _02375_ _02440_ _02441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09937__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10256_ _05012_ memory\[46\]\[3\] _05006_ _05013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_167_3583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12104__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10187_ _04974_ _00159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12449__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14995_ _02034_ clknet_leaf_68_clk_i memory\[38\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12544__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13946_ _00985_ clknet_leaf_388_clk_i memory\[8\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09413__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xload_slew75 _03452_ net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_18_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06923__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13877_ _00916_ clknet_leaf_66_clk_i memory\[39\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15616_ _00575_ clknet_leaf_326_clk_i memory\[58\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12828_ _06603_ _02223_ _02225_ _02227_ _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_16_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15547_ _00506_ clknet_leaf_378_clk_i memory\[55\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12759_ _06467_ _02152_ _02159_ _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_16_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_182_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15478_ _00437_ clknet_leaf_266_clk_i memory\[53\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14429_ _01468_ clknet_leaf_360_clk_i memory\[21\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08428__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09970_ _04639_ memory\[41\]\[31\] _04824_ _04859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08699__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08921_ _04185_ memory\[27\]\[1\] _04286_ _04288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12688__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08852_ _04251_ _01627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08498__I _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08600__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07803_ _03662_ _01167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08783_ _04203_ memory\[25\]\[10\] _04204_ _04205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07734_ _03187_ memory\[63\]\[20\] _03625_ _03626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_88_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09323__S _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07665_ _03566_ _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_49_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13353__B _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09404_ _04543_ _01887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07596_ _03529_ _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_48_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12299__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09122__I _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09335_ _04191_ memory\[33\]\[4\] _04502_ _04507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10474__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09266_ _04470_ _01822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_124_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08217_ _03899_ _01344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09197_ _04189_ memory\[31\]\[3\] _04430_ _04434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10226__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08148_ _03762_ memory\[29\]\[5\] _03857_ _03863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09092__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12471__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08079_ _03825_ _01280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10110_ _04573_ memory\[44\]\[0\] _04933_ _04934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08402__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11090_ _05068_ memory\[57\]\[30\] _05434_ _05468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12679__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12432__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11827__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10041_ _04896_ _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_145_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13800_ _00839_ clknet_leaf_208_clk_i memory\[16\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_49_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11992_ memory\[22\]\[6\] memory\[23\]\[6\] _06062_ _06202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14780_ _01819_ clknet_leaf_427_clk_i memory\[32\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09233__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13731_ _03074_ _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_123_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10943_ _05390_ _00499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10379__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12851__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11562__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13662_ memory\[44\]\[31\] memory\[45\]\[31\] _05678_ _03049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10874_ _05353_ _00467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15401_ _00360_ clknet_leaf_292_clk_i memory\[51\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12613_ _06813_ _06814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_151_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13593_ _02980_ _02981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12603__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12454__I1 memory\[39\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07688__S _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12544_ memory\[24\]\[14\] memory\[25\]\[14\] memory\[26\]\[14\] memory\[27\]\[14\]
+ _06472_ _06611_ _06746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08871__I _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15332_ _00291_ clknet_leaf_282_clk_i memory\[4\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12475_ _06677_ _06678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15263_ _00222_ clknet_leaf_417_clk_i memory\[47\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_401_clk_i clknet_5_3__leaf_clk_i clknet_leaf_401_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10217__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14214_ _01253_ clknet_leaf_201_clk_i memory\[12\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11426_ _05646_ _00726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15194_ _00153_ clknet_leaf_445_clk_i memory\[44\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14145_ _01184_ clknet_leaf_308_clk_i memory\[7\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11357_ memory\[61\]\[27\] _03208_ _05602_ _05610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10308_ _05005_ _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_416_clk_i clknet_5_2__leaf_clk_i clknet_leaf_416_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14076_ _01115_ clknet_leaf_311_clk_i memory\[63\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_326_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11288_ _03365_ memory\[60\]\[27\] _05565_ _05573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13027_ _02213_ _02423_ _02352_ _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10239_ _05001_ _00184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_182_3867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10940__I1 _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13095__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07149__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14978_ _02017_ clknet_leaf_402_clk_i memory\[38\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13929_ _00968_ clknet_leaf_212_clk_i memory\[8\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08897__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07450_ _03473_ _01003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07381_ _03181_ memory\[8\]\[18\] _03426_ _03435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09120_ _04392_ _01754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10456__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08781__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12517__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09051_ _04247_ memory\[28\]\[31\] _04321_ _04356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_6_Right_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08002_ _03159_ _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_167_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11848__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08222__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09953_ _04850_ _00049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08904_ _04278_ _01652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12756__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07388__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09884_ _04621_ memory\[40\]\[22\] _04811_ _04814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08835_ _04239_ memory\[25\]\[27\] _04225_ _04240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10931__I1 _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12508__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_50_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08766_ _03140_ _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_68_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input11_I data_i[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07717_ _03163_ memory\[63\]\[12\] _03614_ _03617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10199__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08888__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08697_ _03766_ memory\[24\]\[7\] _04146_ _04154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_140_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09988__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10695__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07648_ _03580_ _01094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_64_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07579_ _03543_ _01062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_81_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10927__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10447__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09318_ _04497_ _01847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12061__A2 _06239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10590_ _05202_ _00334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_275_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07301__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09249_ _04241_ memory\[31\]\[28\] _04452_ _04461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13102__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12260_ _06445_ _06457_ _06465_ _06466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09065__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07100__I _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11211_ _05532_ _00625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09765__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12191_ memory\[24\]\[9\] memory\[25\]\[9\] memory\[26\]\[9\] memory\[27\]\[9\] _05778_
+ _05922_ _06398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_5_7__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09228__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11142_ _03355_ memory\[58\]\[22\] _05493_ _05496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput43 net43 data_o[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08132__S _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput54 net54 data_o[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_9_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11557__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput65 net65 data_o[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11073_ _05459_ _00560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07379__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10024_ _04625_ memory\[42\]\[24\] _04883_ _04888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14901_ _01940_ clknet_leaf_74_clk_i memory\[35\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14832_ _01871_ clknet_leaf_77_clk_i memory\[33\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12419__A4 _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14763_ _01802_ clknet_leaf_130_clk_i memory\[31\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11975_ _05753_ _06184_ _05757_ _06185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__09898__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13714_ _03088_ _00774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__15495__CLK clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10926_ _05381_ _00491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14694_ _01733_ clknet_leaf_252_clk_i memory\[2\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10837__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13645_ _05759_ _03031_ _03032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10857_ _05344_ _00459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_186_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08307__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_340_clk_i clknet_5_8__leaf_clk_i clknet_leaf_340_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_54_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13576_ _03450_ _02956_ _02963_ _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_10788_ _05039_ memory\[53\]\[16\] _05301_ _05308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_59_Right_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15315_ _00274_ clknet_leaf_158_clk_i memory\[48\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12527_ memory\[38\]\[14\] memory\[39\]\[14\] _06728_ _06729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13001__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15246_ _00205_ clknet_leaf_272_clk_i memory\[46\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12458_ _06446_ _06656_ _06658_ _06660_ _06661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_23_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11668__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11409_ _05637_ _00718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_355_clk_i clknet_5_2__leaf_clk_i clknet_leaf_355_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15177_ _00136_ clknet_leaf_32_clk_i memory\[44\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12389_ _06446_ _06588_ _06590_ _06592_ _06593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_111_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10610__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14128_ _01167_ clknet_leaf_120_clk_i memory\[6\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06950_ net12 _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14059_ _01098_ clknet_leaf_209_clk_i memory\[10\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08977__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_68_Right_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_input3_I address_i[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06881_ _03112_ _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_4
XFILLER_0_101_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10913__I1 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08620_ _04113_ _01533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08551_ _04076_ _01501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07502_ memory\[59\]\[8\] _03325_ _03493_ _03502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08482_ _03756_ memory\[21\]\[2\] _04037_ _04040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12291__A2 _06495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07433_ _03464_ _00995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10747__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13123__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_77_Right_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07364_ _03414_ _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_130_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_308_clk_i clknet_5_14__leaf_clk_i clknet_leaf_308_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09103_ _04231_ memory\[2\]\[23\] _04380_ _04384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07295_ _03389_ _00932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09034_ _04347_ _01713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09047__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06960__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12426__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10482__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_57_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_86_Right_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09936_ _04841_ _00041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07791__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__A2 _06036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09867_ _04604_ memory\[40\]\[14\] _04800_ _04805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_142_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12710__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10904__I1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08818_ _04228_ _01616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09770__I1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09798_ _04767_ _02057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07781__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08749_ _03110_ _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_120_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11760_ memory\[44\]\[3\] memory\[45\]\[3\] _05749_ _05973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_96_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10711_ _05267_ _00390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_95_Right_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_166_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11691_ memory\[44\]\[2\] memory\[45\]\[2\] _05749_ _05905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11880__I2 memory\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_166_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13430_ _02375_ _02820_ _02821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_14_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10642_ memory\[51\]\[11\] _03159_ _05229_ _05231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06934__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09286__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13361_ _02494_ _02748_ _02750_ _02752_ _02753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10573_ _05029_ memory\[50\]\[11\] _05192_ _05194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_118_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11793__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15100_ _00059_ clknet_leaf_440_clk_i memory\[42\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_118_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12312_ memory\[14\]\[11\] memory\[15\]\[11\] _06302_ _06517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13292_ memory\[28\]\[25\] memory\[29\]\[25\] _02495_ _02685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15031_ _02070_ clknet_leaf_56_clk_i memory\[3\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12243_ _06448_ _06449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10392__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12174_ memory\[38\]\[9\] memory\[39\]\[9\] _06039_ _06381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_2_Left_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11125_ _03338_ memory\[58\]\[14\] _05482_ _05487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13298__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11056_ _05450_ _00552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13208__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10007_ _04608_ memory\[42\]\[16\] _04872_ _04879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12112__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07772__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14815_ _01854_ clknet_leaf_424_clk_i memory\[33\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15795_ _00754_ clknet_leaf_88_clk_i net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14746_ _01785_ clknet_leaf_26_clk_i memory\[30\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11958_ memory\[14\]\[6\] memory\[15\]\[6\] _05720_ _06168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_177_3777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_177_3788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10909_ _05372_ _00483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14677_ _01716_ clknet_leaf_83_clk_i memory\[28\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11889_ _06024_ _06095_ _06097_ _06099_ _06100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_172_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13628_ _05705_ _03014_ _05756_ _03015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08037__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11084__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10366__I _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13559_ _02902_ _02917_ _02932_ _02947_ _02948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__07876__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10831__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07080_ _03200_ memory\[16\]\[24\] _03251_ _03256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09029__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12408__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_294_clk_i clknet_5_14__leaf_clk_i clknet_leaf_294_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15229_ _00188_ clknet_leaf_418_clk_i memory\[46\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07982_ _03761_ _01247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13289__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_223_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09721_ _04726_ _02021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06933_ net8 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09201__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13384__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09652_ _04595_ memory\[37\]\[10\] _04689_ _04690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_232_clk_i clknet_5_26__leaf_clk_i clknet_leaf_232_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_179_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_18__f_clk_i clknet_2_2_0_clk_i clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_171_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08603_ _04103_ _01526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09583_ _04641_ _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_26_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08534_ _03808_ memory\[21\]\[27\] _04059_ _04067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_26_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13461__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11311__I1 _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09331__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08465_ _04030_ _01461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_247_clk_i clknet_5_26__leaf_clk_i clknet_leaf_247_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07416_ memory\[49\]\[0\] _03303_ _03455_ _03456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_46_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13213__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08396_ _03806_ memory\[1\]\[26\] _03987_ _03994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07347_ _03417_ _00956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10276__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07278_ memory\[11\]\[1\] _03311_ _03379_ _03381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09017_ _04338_ _01705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_13_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_113_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10940__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09919_ _04832_ _00033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08410__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12440__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12930_ memory\[12\]\[20\] memory\[13\]\[20\] _06714_ _02328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06929__I net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output42_I net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07754__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12861_ _06851_ _02259_ _02260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14600_ _01639_ clknet_leaf_180_clk_i memory\[26\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11812_ _05675_ _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_159_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15580_ _00539_ clknet_leaf_328_clk_i memory\[57\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12792_ _02191_ _02192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_159_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_425_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09241__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14531_ _01570_ clknet_leaf_355_clk_i memory\[24\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11743_ _05710_ _05955_ _05956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12666__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13204__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09259__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14462_ _01501_ clknet_leaf_352_clk_i memory\[22\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11674_ _05700_ _05883_ _05885_ _05887_ _05888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_166_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13698__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13413_ _02213_ _02803_ _02352_ _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_148_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10625_ memory\[51\]\[3\] _03134_ _05218_ _05222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14393_ _01432_ clknet_leaf_54_clk_i memory\[1\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_172_3685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11766__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07696__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_172_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10813__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10556_ _05012_ memory\[50\]\[3\] _05181_ _05185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13344_ memory\[32\]\[26\] memory\[33\]\[26\] memory\[34\]\[26\] memory\[35\]\[26\]
+ _02205_ _02345_ _02736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_109_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12615__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_133_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13275_ _05768_ _02663_ _02665_ _02667_ _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10487_ _05148_ _00285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15014_ _02053_ clknet_leaf_252_clk_i memory\[3\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12226_ memory\[6\]\[10\] memory\[7\]\[10\] _06431_ _06432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_184_Right_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12157_ memory\[4\]\[9\] memory\[5\]\[9\] _06156_ _06364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10850__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07993__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11108_ _03321_ memory\[58\]\[6\] _05471_ _05478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09416__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08320__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13366__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12088_ _06159_ _06295_ _06018_ _06296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13446__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11039_ _05441_ _00544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_179_3817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12777__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_97_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15778_ _00737_ clknet_leaf_337_clk_i net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__09498__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_115_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14729_ _01768_ clknet_leaf_132_clk_i memory\[30\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08250_ _03796_ memory\[17\]\[21\] _03915_ _03917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07201_ memory\[39\]\[9\] _03327_ _03309_ _03328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11057__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08181_ _03880_ _01327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07132_ _03172_ memory\[13\]\[15\] _03279_ _03285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_31_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09670__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Left_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07063_ _03175_ memory\[16\]\[16\] _03240_ _03247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09422__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12182__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_151_Right_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_374_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07984__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07965_ _03748_ _03264_ _03123_ _03749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_96_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_171_clk_i clknet_5_30__leaf_clk_i clknet_leaf_171_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09704_ _04717_ _02013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06916_ _03142_ _00800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07736__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07896_ _03111_ memory\[19\]\[0\] _03711_ _03712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13682__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_74_Left_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09635_ _04579_ memory\[37\]\[2\] _04678_ _04681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11591__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09566_ _04644_ _01948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_186_clk_i clknet_5_29__leaf_clk_i clknet_leaf_186_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09061__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08517_ _03791_ memory\[21\]\[19\] _04048_ _04058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11296__I0 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09497_ _03159_ _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08161__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11996__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08448_ _04021_ _01453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08379_ _03789_ memory\[1\]\[18\] _03976_ _03985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11748__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10410_ _05070_ memory\[47\]\[31\] _05072_ _05107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_78_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Left_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11390_ _03329_ memory\[62\]\[10\] _05627_ _05628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_115_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_150_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10341_ _03220_ _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_131_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_124_clk_i clknet_5_23__leaf_clk_i clknet_leaf_124_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_182_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13060_ memory\[54\]\[22\] memory\[55\]\[22\] _02312_ _02456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_111_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10272_ _05023_ _00195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09413__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13596__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12011_ _06146_ _06219_ _05687_ _06220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11220__I0 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11920__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07975__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08140__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_139_clk_i clknet_5_22__leaf_clk_i clknet_leaf_139_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_92_Left_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_119_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13962_ _01001_ clknet_leaf_238_clk_i memory\[49\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07727__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13673__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15701_ _00660_ clknet_leaf_161_clk_i memory\[60\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12913_ _02310_ _02311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12597__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13893_ _00932_ clknet_leaf_298_clk_i memory\[11\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15632_ _00591_ clknet_leaf_178_clk_i memory\[58\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12844_ _02167_ _02242_ _06690_ _02243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_17_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15563_ _00522_ clknet_leaf_231_clk_i memory\[56\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_174_3725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12775_ memory\[52\]\[18\] memory\[53\]\[18\] _06832_ _02175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08152__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11006__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14514_ _01553_ clknet_leaf_101_clk_i memory\[23\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11726_ _05660_ _05938_ _05665_ _05939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_138_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15494_ _00453_ clknet_leaf_287_clk_i memory\[54\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14445_ _01484_ clknet_leaf_188_clk_i memory\[21\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11657_ memory\[56\]\[2\] memory\[57\]\[2\] memory\[58\]\[2\] memory\[59\]\[2\] _05670_
+ _05671_ _05871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_36_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13221__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10608_ _05064_ memory\[50\]\[28\] _05203_ _05212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14376_ _01415_ clknet_leaf_249_clk_i memory\[1\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09652__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11588_ _05803_ _00731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13327_ memory\[6\]\[26\] memory\[7\]\[26\] _02322_ _02719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10539_ _05175_ _00310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13036__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13258_ memory\[48\]\[25\] memory\[49\]\[25\] memory\[50\]\[25\] memory\[51\]\[25\]
+ _05725_ _06839_ _02651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_27_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12209_ _06276_ _06414_ _06001_ _06415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13189_ _02170_ _02582_ _02583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_86_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11911__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09146__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13176__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12080__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07750_ _03212_ memory\[63\]\[28\] _03625_ _03634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07681_ _03597_ _01110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09420_ _04208_ memory\[34\]\[12\] _04549_ _04552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07894__A2 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13416__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11278__I0 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09351_ _04515_ _01862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11978__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08302_ _03944_ _01384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09282_ _04206_ memory\[32\]\[11\] _04477_ _04479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_185_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08233_ _03779_ memory\[17\]\[13\] _03904_ _03908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10755__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08164_ _03871_ _01319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_95_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_41_clk_i clknet_5_7__leaf_clk_i clknet_leaf_41_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09643__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07115_ _03147_ memory\[13\]\[7\] _03268_ _03276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08095_ _03779_ memory\[15\]\[13\] _03830_ _03834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07046_ _03150_ memory\[16\]\[8\] _03229_ _03238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_73_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_73_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12155__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_56_clk_i clknet_5_19__leaf_clk_i clknet_leaf_56_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10490__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08997_ _04193_ memory\[28\]\[5\] _04322_ _04328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_120_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07948_ _03203_ memory\[19\]\[25\] _03733_ _03739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08895__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07879_ _03702_ _01203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_3_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09618_ _04671_ _01973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10890_ _05361_ _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_156_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11269__I0 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09549_ _03211_ _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_104_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_4047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13105__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12560_ _06760_ _06761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09882__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11511_ memory\[8\]\[0\] memory\[9\]\[0\] memory\[10\]\[0\] memory\[11\]\[0\] _05725_
+ _05726_ _05727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_65_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10492__I1 memory\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10665__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12491_ _06279_ _06692_ _06693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_149_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13266__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13041__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14230_ _01269_ clknet_leaf_110_clk_i memory\[12\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11442_ _05657_ _05658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06942__I net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12394__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_45_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14161_ _01200_ clknet_leaf_119_clk_i memory\[7\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11373_ _03313_ memory\[62\]\[2\] _05616_ _05619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12880__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_46_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13112_ memory\[22\]\[22\] memory\[23\]\[22\] _06751_ _02508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10324_ _05058_ memory\[46\]\[25\] _05048_ _05059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14092_ _01131_ clknet_leaf_224_clk_i memory\[63\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13043_ memory\[16\]\[21\] memory\[17\]\[21\] memory\[18\]\[21\] memory\[19\]\[21\]
+ _02233_ _02376_ _02440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10255_ _03134_ _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_30_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12697__A2 _06862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07948__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10186_ _04583_ memory\[45\]\[4\] _04969_ _04974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_128_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12449__A2 _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13646__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14994_ _02033_ clknet_leaf_68_clk_i memory\[38\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13497__I1 net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13945_ _00984_ clknet_leaf_132_clk_i memory\[8\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08373__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13216__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10180__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13876_ _00915_ clknet_leaf_67_clk_i memory\[39\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15615_ _00574_ clknet_leaf_328_clk_i memory\[58\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12827_ _06610_ _02226_ _02227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_5_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10639__I _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_322_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15546_ _00505_ clknet_leaf_379_clk_i memory\[55\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12758_ _06476_ _02154_ _02156_ _02158_ _02159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08109__I _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09873__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11709_ memory\[24\]\[2\] memory\[25\]\[2\] memory\[26\]\[2\] memory\[27\]\[2\] _05778_
+ _05922_ _05923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_71_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10575__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15477_ _00436_ clknet_leaf_263_clk_i memory\[53\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12689_ memory\[20\]\[16\] memory\[21\]\[16\] _06477_ _02091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14428_ _01467_ clknet_leaf_361_clk_i memory\[21\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09625__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14359_ _01398_ clknet_leaf_107_clk_i memory\[18\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07884__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Left_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12137__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08920_ _04287_ _01659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08851_ _04181_ memory\[26\]\[0\] _04250_ _04251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07802_ _03187_ memory\[6\]\[20\] _03661_ _03662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08782_ _04182_ _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13637__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07733_ _03602_ _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_0_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11933__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07664_ _03588_ _01102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_49_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07124__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_148_Left_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09403_ _04191_ memory\[34\]\[4\] _04538_ _04543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07595_ _03551_ _01070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10549__I _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08116__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12299__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09334_ _04506_ _01854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__I1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12764__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09265_ _04189_ memory\[32\]\[3\] _04466_ _04470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08216_ _03762_ memory\[17\]\[5\] _03893_ _03899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09196_ _04433_ _01789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11423__I0 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08147_ _03862_ _01311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_157_Left_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12471__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08078_ _03762_ memory\[15\]\[5\] _03819_ _03825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12128__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07029_ _03228_ _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_140_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10040_ _03376_ _04787_ _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_8_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_145_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_271_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13628__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12939__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11991_ _06200_ _06201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_106_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_166_Left_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12300__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11734__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13730_ _03096_ _00782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10942_ memory\[55\]\[24\] _03199_ _05385_ _05390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10162__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07034__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13661_ _05654_ _03043_ _03045_ _03047_ _03048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10873_ _05056_ memory\[54\]\[24\] _05348_ _05353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08107__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15400_ _00359_ clknet_leaf_292_clk_i memory\[51\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12612_ memory\[20\]\[15\] memory\[21\]\[15\] _06477_ _06813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07969__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13592_ memory\[36\]\[30\] memory\[37\]\[30\] _05656_ _02980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15331_ _00290_ clknet_leaf_337_clk_i memory\[4\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12543_ _06607_ _06744_ _06195_ _06745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_136_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__I1 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15262_ _00221_ clknet_leaf_416_clk_i memory\[47\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12474_ memory\[20\]\[13\] memory\[21\]\[13\] _06477_ _06677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09607__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14213_ _01252_ clknet_leaf_288_clk_i memory\[12\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11425_ _03365_ memory\[62\]\[27\] _05638_ _05646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15193_ _00152_ clknet_leaf_23_clk_i memory\[44\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07094__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14144_ _01183_ clknet_leaf_308_clk_i memory\[7\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11356_ _05609_ _00693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_186_3960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10307_ _03186_ _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12115__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14075_ _01114_ clknet_leaf_386_clk_i memory\[10\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11287_ _05572_ _00661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13026_ memory\[46\]\[21\] memory\[47\]\[21\] _06596_ _02423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10238_ _04635_ memory\[45\]\[29\] _04991_ _05001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08594__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10169_ _04964_ _00151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13619__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07008__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09424__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13454__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14977_ _02016_ clknet_leaf_421_clk_i memory\[38\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08346__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13928_ _00967_ clknet_leaf_212_clk_i memory\[8\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13859_ _00898_ clknet_leaf_402_clk_i memory\[39\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07380_ _03434_ _00972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09846__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15529_ _00488_ clknet_leaf_290_clk_i memory\[55\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09050_ _04355_ _01721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12358__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08001_ _03774_ _01253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08503__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11928__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12025__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09952_ _04621_ memory\[41\]\[22\] _04847_ _04850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08903_ _04235_ memory\[26\]\[25\] _04272_ _04278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07119__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09883_ _04813_ _00016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08585__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08834_ _03208_ _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_32_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10392__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08765_ _04192_ _01599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_68_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11716__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07716_ _03616_ _01126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08696_ _04153_ _01569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06899__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07647_ _03160_ memory\[10\]\[11\] _03578_ _03580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07789__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07578_ _03160_ memory\[0\]\[11\] _03541_ _03543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_81_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09317_ _04241_ memory\[32\]\[28\] _04488_ _04497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_218_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09462__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12061__A3 _06254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11104__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09248_ _04460_ _01814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09179_ _04239_ memory\[30\]\[27\] _04416_ _04424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09065__I1 memory\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07076__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11210_ _03355_ memory\[5\]\[22\] _05529_ _05532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12190_ _05918_ _06396_ _06195_ _06397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_114_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13539__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11141_ _05495_ _00592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xoutput44 net44 data_o[13] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_147_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput55 net55 data_o[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput66 net66 data_o[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_11072_ _05050_ memory\[57\]\[21\] _05457_ _05459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_164_3532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12521__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10023_ _04887_ _00082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14900_ _01939_ clknet_leaf_74_clk_i memory\[35\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10383__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14831_ _01870_ clknet_leaf_63_clk_i memory\[33\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08328__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11573__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14762_ _01801_ clknet_leaf_131_clk_i memory\[31\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11974_ memory\[46\]\[6\] memory\[47\]\[6\] _05907_ _06184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10135__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_98_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13713_ _03332_ memory\[9\]\[11\] _03086_ _03088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10925_ memory\[55\]\[16\] _03174_ _05374_ _05381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14693_ _01732_ clknet_leaf_360_clk_i memory\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13644_ memory\[0\]\[31\] memory\[1\]\[31\] memory\[2\]\[31\] memory\[3\]\[31\] _05784_
+ _03226_ _03031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_39_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10856_ _05039_ memory\[54\]\[16\] _05337_ _05344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12588__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13575_ _05715_ _02958_ _02960_ _02962_ _02963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_125_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10787_ _05307_ _00426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07303__I1 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15314_ _00273_ clknet_leaf_158_clk_i memory\[48\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12526_ _05661_ _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_41_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15245_ _00204_ clknet_leaf_277_clk_i memory\[46\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12457_ _06453_ _06659_ _06660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_136_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07067__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11408_ _03348_ memory\[62\]\[19\] _05627_ _05637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15176_ _00135_ clknet_leaf_32_clk_i memory\[44\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12388_ _06453_ _06591_ _06592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_184_3908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_184_3919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14127_ _01166_ clknet_leaf_219_clk_i memory\[6\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11339_ _05600_ _00685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14058_ _01097_ clknet_leaf_212_clk_i memory\[10\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08567__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11684__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13009_ memory\[12\]\[21\] memory\[13\]\[21\] _06714_ _02406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06880_ net4 _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09154__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11483__I _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08550_ _03756_ memory\[22\]\[2\] _04073_ _04076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08993__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10126__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11618__A3 _05832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12815__A2 _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12371__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07501_ _03501_ _01026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08481_ _04039_ _01468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10677__I1 _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07542__I1 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07432_ memory\[49\]\[8\] _03325_ _03455_ _03464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07402__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12528__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07363_ _03425_ _00964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09102_ _04383_ _01745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07294_ memory\[11\]\[9\] _03327_ _03379_ _03389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09033_ _04229_ memory\[28\]\[22\] _04344_ _04347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10763__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12426__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09329__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08233__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07758__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12751__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09935_ _04604_ memory\[41\]\[14\] _04836_ _04841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08558__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09866_ _04804_ _00008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_142_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__A3 _06052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08817_ _04227_ memory\[25\]\[21\] _04225_ _04228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11607__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09797_ memory\[3\]\[14\] _03168_ _04762_ _04767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_400_clk_i clknet_5_1__leaf_clk_i clknet_leaf_400_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09999__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08748_ _04180_ _01594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10003__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08679_ memory\[23\]\[31\] _03373_ _04109_ _04144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10938__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10710_ _05029_ memory\[52\]\[11\] _05265_ _05267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11690_ _05732_ _05899_ _05901_ _05903_ _05904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xclkbuf_leaf_415_clk_i clknet_5_2__leaf_clk_i clknet_leaf_415_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10641_ _05230_ _00357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_369_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13360_ _02501_ _02751_ _02752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_146_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10572_ _05193_ _00325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_165_Right_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_118_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12311_ _06515_ _06516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12990__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10673__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13291_ _02336_ _02676_ _02683_ _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_134_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09239__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15030_ _02069_ clknet_leaf_58_clk_i memory\[3\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12242_ memory\[36\]\[10\] memory\[37\]\[10\] _06447_ _06448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06950__I net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11568__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12742__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_421_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12173_ _06379_ _06380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_82_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11124_ _05486_ _00584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11055_ _05033_ memory\[57\]\[13\] _05446_ _05450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10356__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10006_ _04878_ _00074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12399__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14814_ _01853_ clknet_leaf_424_clk_i memory\[33\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15794_ _00753_ clknet_leaf_58_clk_i net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14745_ _01784_ clknet_leaf_60_clk_i memory\[30\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11957_ _06166_ _06167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10848__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11481__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10908_ memory\[55\]\[8\] _03149_ _05363_ _05372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14676_ _01715_ clknet_leaf_94_clk_i memory\[28\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08318__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_177_3789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11888_ _06031_ _06098_ _06099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_103_Left_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13627_ memory\[62\]\[31\] memory\[63\]\[31\] _02448_ _03014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10839_ _05022_ memory\[54\]\[8\] _05326_ _05335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13558_ _02358_ _02939_ _02946_ _02947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_82_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_132_Right_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12981__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12509_ _06162_ _06710_ _06711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10583__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13489_ _02878_ _02879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12408__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_93_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15228_ _00187_ clknet_leaf_421_clk_i memory\[46\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11478__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12733__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15159_ _00118_ clknet_leaf_6_clk_i memory\[43\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__S _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07981_ _03760_ memory\[12\]\[4\] _03752_ _03761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13289__A2 _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09720_ _04595_ memory\[38\]\[10\] _04725_ _04726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06932_ _03154_ _00804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12303__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07691__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09651_ _04677_ _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10898__I1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08602_ _03808_ memory\[22\]\[27\] _04095_ _04103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09582_ _04652_ _01956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12344__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_26_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08533_ _04066_ _01493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08712__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07515__I1 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11472__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08464_ _03806_ memory\[20\]\[26\] _04023_ _04030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07132__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07415_ _03454_ _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_18_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_370_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08395_ _03993_ _01428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07346_ _03129_ memory\[8\]\[1\] _03415_ _03417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11589__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07277_ _03380_ _00923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09016_ _04212_ memory\[28\]\[14\] _04333_ _04338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09059__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_170_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08779__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10292__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09918_ _04587_ memory\[41\]\[6\] _04825_ _04832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12213__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07307__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09849_ _04795_ _00000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12860_ memory\[0\]\[19\] memory\[1\]\[19\] memory\[2\]\[19\] memory\[3\]\[19\] _06709_
+ _06779_ _02259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09522__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11811_ _05700_ _06016_ _06019_ _06022_ _06023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12947__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12791_ memory\[12\]\[18\] memory\[13\]\[18\] _06714_ _02191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_354_clk_i clknet_5_2__leaf_clk_i clknet_leaf_354_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14530_ _01569_ clknet_leaf_409_clk_i memory\[24\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11742_ memory\[0\]\[3\] memory\[1\]\[3\] memory\[2\]\[3\] memory\[3\]\[3\] _05711_
+ _03748_ _05955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_96_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08138__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07042__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14461_ _01500_ clknet_leaf_365_clk_i memory\[22\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11673_ _05710_ _05886_ _05887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13412_ memory\[46\]\[27\] memory\[47\]\[27\] _02487_ _02803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10624_ _05221_ _00349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_12_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14392_ _01431_ clknet_leaf_55_clk_i memory\[1\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_369_clk_i clknet_5_9__leaf_clk_i clknet_leaf_369_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_115_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_172_3686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12682__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13343_ _02341_ _02734_ _05708_ _02735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10555_ _05184_ _00317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13274_ _05777_ _02666_ _02667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_45_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10486_ _05010_ memory\[4\]\[2\] _05145_ _05148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15013_ _02052_ clknet_leaf_339_clk_i memory\[3\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12225_ _05661_ _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10577__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12156_ _05651_ _06355_ _06362_ _06363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_11107_ _05477_ _00576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12123__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12087_ memory\[6\]\[8\] memory\[7\]\[8\] _05706_ _06295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_307_clk_i clknet_5_14__leaf_clk_i clknet_leaf_307_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09195__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11038_ _05016_ memory\[57\]\[5\] _05435_ _05441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08942__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07016__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09432__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12989_ memory\[62\]\[21\] memory\[63\]\[21\] _06557_ _02386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15777_ _00736_ clknet_leaf_344_clk_i net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_111_Left_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14728_ _01767_ clknet_leaf_180_clk_i memory\[30\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14659_ _01698_ clknet_leaf_355_clk_i memory\[28\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07200_ _03152_ _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_129_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08180_ _03793_ memory\[29\]\[20\] _03879_ _03880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07131_ _03284_ _00873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07062_ _03246_ _00842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_120_Left_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12706__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13754__I0 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12557__I1 net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10568__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11001__I _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09607__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_54_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08511__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_317_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11936__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12033__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07964_ _03747_ _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_96_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_71_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09703_ _04579_ memory\[38\]\[2\] _04714_ _04717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13131__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06915_ _03141_ memory\[14\]\[5\] _03126_ _03142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07895_ _03710_ _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08933__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09634_ _04680_ _01980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12767__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09565_ _04577_ memory\[36\]\[1\] _04642_ _04644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10488__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08516_ _04057_ _01485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09496_ _04597_ _01925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08447_ _03789_ memory\[20\]\[18\] _04012_ _04021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13198__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07797__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_154_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_92_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08378_ _03984_ _01420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07329_ _03407_ _00948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12208__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07596__I _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11112__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07672__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10340_ _05069_ _00217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10271_ _05022_ memory\[46\]\[8\] _05006_ _05023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13370__A1 _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12010_ memory\[54\]\[7\] memory\[55\]\[7\] _05684_ _06219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13547__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13039__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09177__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13961_ _01000_ clknet_leaf_295_clk_i memory\[49\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12878__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15700_ _00659_ clknet_leaf_162_clk_i memory\[60\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12912_ memory\[52\]\[20\] memory\[53\]\[20\] _06832_ _02310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_41_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13892_ _00931_ clknet_leaf_299_clk_i memory\[11\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10731__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_293_clk_i clknet_5_15__leaf_clk_i clknet_leaf_293_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12843_ memory\[62\]\[19\] memory\[63\]\[19\] _06557_ _02242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15631_ _00590_ clknet_leaf_243_clk_i memory\[58\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09629__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10398__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11436__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15562_ _00521_ clknet_leaf_231_clk_i memory\[56\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12774_ _02163_ _02166_ _02169_ _02173_ _02174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_185_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14513_ _01552_ clknet_leaf_104_clk_i memory\[23\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11725_ memory\[62\]\[3\] memory\[63\]\[3\] _05868_ _05938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15493_ _00452_ clknet_leaf_313_clk_i memory\[54\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13189__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14444_ _01483_ clknet_leaf_192_clk_i memory\[21\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11656_ _05660_ _05869_ _05665_ _05870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_65_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09101__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12626__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07500__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_266_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12936__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10607_ _05211_ _00342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_182_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14375_ _01414_ clknet_leaf_251_clk_i memory\[1\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11587_ _05801_ net40 _05802_ _05803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11022__S _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13326_ _02717_ _02718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_231_clk_i clknet_5_26__leaf_clk_i clknet_leaf_231_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07663__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10538_ _05062_ memory\[4\]\[27\] _05167_ _05175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13036__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13736__I0 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13257_ _06835_ _02649_ _02178_ _02650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10469_ _05138_ _00277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13361__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12208_ memory\[62\]\[10\] memory\[63\]\[10\] _05868_ _06414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13188_ memory\[56\]\[24\] memory\[57\]\[24\] memory\[58\]\[24\] memory\[59\]\[24\]
+ _06827_ _02171_ _02582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_246_clk_i clknet_5_26__leaf_clk_i clknet_leaf_246_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10660__I _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12139_ _06292_ _06309_ _06330_ _06346_ _06347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_97_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10970__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13113__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08915__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07680_ _03209_ memory\[10\]\[27\] _03589_ _03597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10722__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09162__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15829_ _00788_ clknet_leaf_129_clk_i memory\[9\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09350_ _04206_ memory\[33\]\[11\] _04513_ _04515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08301_ _03779_ memory\[18\]\[13\] _03940_ _03944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09281_ _04478_ _01829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13412__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08232_ _03907_ _01351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08163_ _03777_ memory\[29\]\[12\] _03868_ _03871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07114_ _03275_ _00865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08094_ _03833_ _01287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13727__I0 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11867__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07045_ _03237_ _00834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10771__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09337__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13352__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10570__I _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08996_ _04327_ _01695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13104__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input34_I data_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07947_ _03738_ _01235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12698__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11666__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07878_ _03200_ memory\[7\]\[24\] _03697_ _03702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_3_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09617_ _04629_ memory\[36\]\[26\] _04664_ _04671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12497__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10011__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09548_ _04632_ _01942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_104_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09331__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_4048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07098__A1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12091__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09479_ _04585_ memory\[35\]\[5\] _04575_ _04586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10946__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11510_ _05693_ _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_152_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08416__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12490_ memory\[56\]\[14\] memory\[57\]\[14\] memory\[58\]\[14\] memory\[59\]\[14\]
+ _06138_ _06280_ _06692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_136_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07320__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13266__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12918__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11441_ memory\[60\]\[0\] memory\[61\]\[0\] _05656_ _05657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_61_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14160_ _01199_ clknet_leaf_120_clk_i memory\[7\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07645__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13591__A1 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12394__A2 _06597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11372_ _05618_ _00700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13111_ _02506_ _02507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__11777__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12960__I _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10323_ _03202_ _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_14091_ _01130_ clknet_leaf_225_clk_i memory\[63\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10681__S _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09247__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13042_ _02371_ _02438_ _02373_ _02439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10254_ _05011_ _00189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11576__I _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12697__A3 _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08070__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10185_ _04973_ _00158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07990__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12529__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14993_ _02032_ clknet_leaf_64_clk_i memory\[38\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12401__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13944_ _00983_ clknet_leaf_133_clk_i memory\[8\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_89_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13875_ _00914_ clknet_leaf_61_clk_i memory\[39\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12826_ memory\[24\]\[18\] memory\[25\]\[18\] memory\[26\]\[18\] memory\[27\]\[18\]
+ _06472_ _06611_ _02226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15614_ _00573_ clknet_leaf_326_clk_i memory\[58\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12757_ _06484_ _02157_ _02158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12082__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15545_ _00504_ clknet_leaf_385_clk_i memory\[55\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10856__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11708_ _03747_ _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07884__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15476_ _00435_ clknet_leaf_262_clk_i memory\[53\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12688_ _06603_ _02083_ _02087_ _02089_ _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08326__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14427_ _01466_ clknet_leaf_0_clk_i memory\[20\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_170_clk_i clknet_5_25__leaf_clk_i clknet_leaf_170_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_4_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11639_ _05777_ _05853_ _05854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13582__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07636__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14358_ _01397_ clknet_leaf_107_clk_i memory\[18\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_27__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13309_ _02701_ _00756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14289_ _01328_ clknet_leaf_94_clk_i memory\[29\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_90_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09389__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07964__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_185_clk_i clknet_5_29__leaf_clk_i clknet_leaf_185_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13187__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08061__S _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11486__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08850_ _04249_ _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08061__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11896__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07801_ _03638_ _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08781_ _03155_ _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07732_ _03624_ _01134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11648__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07663_ _03184_ memory\[10\]\[19\] _03578_ _03588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_49_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09402_ _04542_ _01886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_123_clk_i clknet_5_23__leaf_clk_i clknet_leaf_123_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_49_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12110__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07594_ _03184_ memory\[0\]\[19\] _03541_ _03551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07204__I _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09313__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09333_ _04189_ memory\[33\]\[3\] _04502_ _04506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13650__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09264_ _04469_ _01821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07140__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_138_clk_i clknet_5_22__leaf_clk_i clknet_leaf_138_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08215_ _03898_ _01343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09195_ _04187_ memory\[31\]\[2\] _04430_ _04433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_9_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08146_ _03760_ memory\[29\]\[4\] _03857_ _03862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08077_ _03824_ _01279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09067__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07028_ _03225_ _03227_ _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__11187__I0 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08052__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_214_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08979_ _04243_ memory\[27\]\[29\] _04308_ _04318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_145_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13317__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11639__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11990_ memory\[20\]\[6\] memory\[21\]\[6\] _05785_ _06200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07315__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11734__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10941_ _05389_ _00498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13660_ _05668_ _03046_ _03047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10872_ _05352_ _00466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_151_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12611_ _06603_ _06807_ _06809_ _06811_ _06812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_17_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13591_ _03114_ _02971_ _02978_ _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_94_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15330_ _00289_ clknet_leaf_337_clk_i memory\[4\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12542_ memory\[30\]\[14\] memory\[31\]\[14\] _06193_ _06744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08146__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11811__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15261_ _00220_ clknet_leaf_418_clk_i memory\[47\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12473_ _06603_ _06671_ _06673_ _06675_ _06676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_164_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14212_ _01251_ clknet_leaf_276_clk_i memory\[12\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11424_ _05645_ _00725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12998__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15192_ _00151_ clknet_leaf_23_clk_i memory\[44\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14143_ _01182_ clknet_leaf_285_clk_i memory\[7\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_104_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_169_3636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11355_ memory\[61\]\[26\] _03205_ _05602_ _05609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13316__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10306_ _05046_ _00206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_186_3950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14074_ _01113_ clknet_leaf_386_clk_i memory\[10\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11286_ _03363_ memory\[60\]\[26\] _05565_ _05572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11178__I0 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13025_ _02421_ _02422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08043__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11878__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10237_ _05000_ _00183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_182_3869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09705__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10168_ _04633_ memory\[44\]\[28\] _04955_ _04964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14976_ _02015_ clknet_leaf_420_clk_i memory\[38\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10099_ _04927_ _00118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_40_clk_i clknet_5_18__leaf_clk_i clknet_leaf_40_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13927_ _00966_ clknet_leaf_225_clk_i memory\[8\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_0_0_clk_i clknet_0_clk_i clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_88_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_179_Right_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_187_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13858_ _00897_ clknet_leaf_403_clk_i memory\[39\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_416_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_130_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12809_ _05675_ _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_29_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11102__I0 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_55_clk_i clknet_5_19__leaf_clk_i clknet_leaf_55_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13789_ _00828_ clknet_leaf_366_clk_i memory\[16\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07857__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11802__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15528_ _00487_ clknet_leaf_290_clk_i memory\[55\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07482__A1 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15459_ _00418_ clknet_leaf_315_clk_i memory\[53\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08000_ _03772_ memory\[12\]\[10\] _03773_ _03774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_163_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07609__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08282__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11210__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13307__A1 _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09951_ _04849_ _00048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_111_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08902_ _04277_ _01651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08034__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09882_ _04619_ memory\[40\]\[21\] _04811_ _04813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_5_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09615__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08833_ _04238_ _01621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08764_ _04191_ memory\[25\]\[4\] _04183_ _04192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07715_ _03160_ memory\[63\]\[11\] _03614_ _03616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11716__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12294__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08695_ _03764_ memory\[24\]\[6\] _04146_ _04153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_88_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07646_ _03579_ _01093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_140_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_146_Right_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_95_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09350__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_101_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07577_ _03542_ _01061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10496__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07869__I _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09316_ _04496_ _01846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_24_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09462__A2 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12061__A4 _06269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09247_ _04239_ memory\[31\]\[27\] _04452_ _04460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10295__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09178_ _04423_ _01781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_5_9__f_clk_i clknet_2_1_0_clk_i clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_47_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08129_ _03851_ _01304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12216__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11140_ _03353_ memory\[58\]\[21\] _05493_ _05495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_147_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput45 net45 data_o[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput56 net56 data_o[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
Xoutput67 net67 data_o[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_11071_ _05458_ _00559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_164_3533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_365_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12521__A2 _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10022_ _04623_ memory\[42\]\[23\] _04883_ _04887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14830_ _01869_ clknet_leaf_63_clk_i memory\[33\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12886__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14761_ _01800_ clknet_leaf_132_clk_i memory\[31\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11973_ _06182_ _06183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_118_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13712_ _03087_ _00773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10924_ _05380_ _00490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14692_ _01731_ clknet_leaf_377_clk_i memory\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_113_Right_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12037__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13290__B _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13643_ _05752_ _03029_ _05791_ _03030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10855_ _05343_ _00458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__I1 _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13574_ _05724_ _02961_ _02962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_67_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10786_ _05037_ memory\[53\]\[15\] _05301_ _05307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12525_ _06726_ _06727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15313_ _00272_ clknet_leaf_261_clk_i memory\[48\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09994__I _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15244_ _00203_ clknet_leaf_273_clk_i memory\[46\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12456_ memory\[32\]\[13\] memory\[33\]\[13\] memory\[34\]\[13\] memory\[35\]\[13\]
+ _06314_ _06454_ _06659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08604__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13001__A3 _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11407_ _05636_ _00717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08264__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15175_ _00134_ clknet_leaf_31_clk_i memory\[44\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10933__I _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12387_ memory\[32\]\[12\] memory\[33\]\[12\] memory\[34\]\[12\] memory\[35\]\[12\]
+ _06314_ _06454_ _06591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_22_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11030__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14126_ _01165_ clknet_leaf_219_clk_i memory\[6\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10071__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11338_ memory\[61\]\[18\] _03180_ _05591_ _05600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12760__A2 _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14057_ _01096_ clknet_leaf_212_clk_i memory\[10\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11269_ _03346_ memory\[60\]\[18\] _05554_ _05563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07019__I net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13008_ _06844_ _02400_ _02402_ _02404_ _02405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__13560__I1 net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09516__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_85_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14959_ _01998_ clknet_leaf_65_clk_i memory\[37\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07500_ memory\[59\]\[7\] _03323_ _03493_ _03501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12371__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08480_ _03754_ memory\[21\]\[1\] _04037_ _04039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07431_ _03463_ _00994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12028__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_185_Left_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07362_ _03153_ memory\[8\]\[9\] _03415_ _03425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09101_ _04229_ memory\[2\]\[22\] _04380_ _04383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_21_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07293_ _03388_ _00931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13420__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09032_ _04346_ _01712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13528__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11939__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12200__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10843__I _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11875__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09934_ _04840_ _00040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09345__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09755__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09865_ _04602_ memory\[40\]\[13\] _04800_ _04804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_142_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11857__A4 _06068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08816_ _03190_ _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09796_ _04766_ _02056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09507__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08747_ _03816_ memory\[24\]\[31\] _04145_ _04180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08678_ _04143_ _01561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09080__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07629_ _03570_ _01085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12019__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10640_ memory\[51\]\[10\] _03155_ _05229_ _05230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_157_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07297__I1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08494__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10954__S _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10571_ _05026_ memory\[50\]\[10\] _05192_ _05193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12310_ memory\[12\]\[11\] memory\[13\]\[11\] _06025_ _06515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13519__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13290_ _02209_ _02678_ _02680_ _02682_ _02683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_107_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_118_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08424__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12241_ _05655_ _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_32_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12742__A2 _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12172_ memory\[36\]\[9\] memory\[37\]\[9\] _05733_ _06379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10753__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11123_ _03336_ memory\[58\]\[13\] _05482_ _05486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09255__S _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11054_ _05449_ _00551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12050__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10005_ _04606_ memory\[42\]\[15\] _04872_ _04878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_111_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09054__I _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14813_ _01852_ clknet_leaf_428_clk_i memory\[33\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12258__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15793_ _00752_ clknet_leaf_88_clk_i net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14744_ _01783_ clknet_leaf_60_clk_i memory\[30\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11956_ memory\[12\]\[6\] memory\[13\]\[6\] _06025_ _06166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10907_ _05371_ _00482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_177_3779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14675_ _01714_ clknet_leaf_83_clk_i memory\[28\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11887_ memory\[8\]\[5\] memory\[9\]\[5\] memory\[10\]\[5\] memory\[11\]\[5\] _05893_
+ _06032_ _06098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_73_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10838_ _05334_ _00450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13626_ _03012_ _03013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_183_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_41_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07288__I1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13557_ _02367_ _02941_ _02943_ _02945_ _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__11864__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10769_ _05020_ memory\[53\]\[7\] _05290_ _05298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12508_ memory\[0\]\[14\] memory\[1\]\[14\] memory\[2\]\[14\] memory\[3\]\[14\] _06709_
+ _06090_ _06710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_70_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08334__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13488_ memory\[20\]\[28\] memory\[21\]\[28\] _02368_ _02878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_36_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_415 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08237__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12439_ memory\[6\]\[13\] memory\[7\]\[13\] _06431_ _06642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15227_ _00186_ clknet_leaf_0_clk_i memory\[45\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10044__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15158_ _00117_ clknet_leaf_6_clk_i memory\[43\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_39_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14109_ _01148_ clknet_leaf_286_clk_i memory\[6\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07980_ _03137_ _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15089_ _00048_ clknet_leaf_16_clk_i memory\[41\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07460__I1 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09165__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06931_ _03153_ memory\[14\]\[9\] _03126_ _03154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11494__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09650_ _04688_ _01988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10104__S _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08601_ _04102_ _01525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09581_ _04593_ memory\[36\]\[9\] _04642_ _04652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08532_ _03806_ memory\[21\]\[26\] _04059_ _04066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12344__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08509__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08463_ _04029_ _01460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_313_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07414_ _03453_ _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_174_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08394_ _03804_ memory\[1\]\[25\] _03987_ _03993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13213__A3 _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07345_ _03416_ _00955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_72_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_27__f_clk_i clknet_2_3_0_clk_i clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07276_ memory\[11\]\[0\] _03303_ _03379_ _03380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09015_ _04337_ _01704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_131_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09976__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12280__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07451__I1 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09917_ _04831_ _00032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08400__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09848_ _04585_ memory\[40\]\[5\] _04789_ _04795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09803__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09779_ _04757_ _02048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13325__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11810_ _05710_ _06021_ _06022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12790_ _06844_ _02185_ _02187_ _02189_ _02190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_159_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09900__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11741_ _05705_ _05953_ _05708_ _05954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12660__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11672_ memory\[0\]\[2\] memory\[1\]\[2\] memory\[2\]\[2\] memory\[3\]\[2\] _05711_
+ _03748_ _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_14460_ _01499_ clknet_leaf_362_clk_i memory\[22\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_165_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10623_ memory\[51\]\[2\] _03131_ _05218_ _05221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13411_ _02801_ _02802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14391_ _01430_ clknet_leaf_56_clk_i memory\[1\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_12_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13060__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_172_3687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10274__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13342_ memory\[38\]\[26\] memory\[39\]\[26\] _05662_ _02734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10554_ _05010_ memory\[50\]\[2\] _05181_ _05184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08154__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11579__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13273_ memory\[8\]\[25\] memory\[9\]\[25\] memory\[10\]\[25\] memory\[11\]\[25\]
+ _02473_ _05779_ _02666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_133_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10485_ _05147_ _00284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07993__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12224_ _06429_ _06430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15012_ _02051_ clknet_leaf_370_clk_i memory\[3\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_161_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_103_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12155_ _06142_ _06357_ _06359_ _06361_ _06362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12404__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11106_ _03319_ memory\[58\]\[5\] _05471_ _05477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12086_ _06293_ _06294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_34_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11037_ _05440_ _00543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_262_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09713__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15776_ _00735_ clknet_leaf_344_clk_i net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12988_ _02384_ _02385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09512__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14727_ _01766_ clknet_leaf_132_clk_i memory\[30\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11939_ _05689_ _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_115_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14658_ _01697_ clknet_leaf_359_clk_i memory\[28\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08458__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13609_ memory\[30\]\[30\] memory\[31\]\[30\] _05737_ _02997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10594__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11837__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14589_ _01628_ clknet_leaf_406_clk_i memory\[26\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07130_ _03169_ memory\[13\]\[14\] _03279_ _03284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10265__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08064__S _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07130__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11489__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07061_ _03172_ memory\[16\]\[15\] _03240_ _03246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09958__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_54_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07408__S _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_414_clk_i clknet_5_2__leaf_clk_i clknet_leaf_414_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07963_ net2 _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XTAP_TAPCELL_ROW_71_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_71_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09702_ _04716_ _02012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06914_ _03140_ _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07894_ _03225_ _03376_ _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__07207__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09623__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09633_ _04577_ memory\[37\]\[1\] _04678_ _04680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10769__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06944__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13145__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11952__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_429_clk_i clknet_5_1__leaf_clk_i clknet_leaf_429_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09564_ _04643_ _01947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08239__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07143__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08515_ _03789_ memory\[21\]\[18\] _04048_ _04057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08697__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12642__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09495_ _04595_ memory\[35\]\[10\] _04596_ _04597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13690__I0 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08446_ _04020_ _01452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_137_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08449__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08377_ _03787_ memory\[1\]\[17\] _03976_ _03984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11901__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_154_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12245__I1 memory\[39\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10256__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07328_ memory\[11\]\[25\] _03361_ _03401_ _03407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07259_ _03211_ _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_143_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10009__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10270_ _03149_ _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_44_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13370__A2 _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07424__I1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07318__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12005__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13960_ _00999_ clknet_leaf_239_clk_i memory\[49\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12911_ _02163_ _02304_ _02306_ _02308_ _02309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10679__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13891_ _00930_ clknet_leaf_301_clk_i memory\[11\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15630_ _00589_ clknet_leaf_247_clk_i memory\[58\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12842_ _02240_ _02241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07053__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09629__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_17_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11436__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_90_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15561_ _00520_ clknet_leaf_233_clk_i memory\[56\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12773_ _02170_ _02172_ _02173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_174_3716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_68_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14512_ _01551_ clknet_leaf_101_clk_i memory\[23\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_174_3727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11724_ _05936_ _05937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15492_ _00451_ clknet_leaf_313_clk_i memory\[54\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07360__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14443_ _01482_ clknet_leaf_191_clk_i memory\[21\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11655_ memory\[62\]\[2\] memory\[63\]\[2\] _05868_ _05869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_209_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11303__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10247__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10606_ _05062_ memory\[50\]\[27\] _05203_ _05211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14374_ _01413_ clknet_leaf_250_clk_i memory\[1\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11586_ _03122_ _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_51_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_17__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13325_ memory\[4\]\[26\] memory\[5\]\[26\] _05789_ _02717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10537_ _05174_ _00309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10468_ _05060_ memory\[48\]\[26\] _05131_ _05138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13256_ memory\[54\]\[25\] memory\[55\]\[25\] _02312_ _02649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12207_ _06412_ _06413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13187_ _02167_ _02580_ _05756_ _02581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10399_ _05101_ _00244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12138_ _05767_ _06337_ _06345_ _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_62_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12069_ memory\[62\]\[8\] memory\[63\]\[8\] _05868_ _06277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09443__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10589__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15828_ _00787_ clknet_leaf_128_clk_i memory\[9\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_56_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15759_ _00718_ clknet_leaf_246_clk_i memory\[62\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08300_ _03943_ _01383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10486__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07898__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09280_ _04203_ memory\[32\]\[10\] _04477_ _04478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08231_ _03777_ memory\[17\]\[12\] _03904_ _03907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10238__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08162_ _03870_ _01318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07103__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07113_ _03144_ memory\[13\]\[6\] _03268_ _03275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08093_ _03777_ memory\[15\]\[12\] _03830_ _03833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08851__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07044_ _03147_ memory\[16\]\[7\] _03229_ _03237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08522__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12235__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_73_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13352__A2 _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_353_clk_i clknet_5_2__leaf_clk_i clknet_leaf_353_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_41_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07138__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10410__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08995_ _04191_ memory\[28\]\[4\] _04322_ _04327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11883__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06977__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07946_ _03200_ memory\[19\]\[24\] _03733_ _03738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_368_clk_i clknet_5_9__leaf_clk_i clknet_leaf_368_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_input27_I data_i[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_5_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13383__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07877_ _03701_ _01202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12778__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_158_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09616_ _04670_ _01972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07590__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10298__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12615__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09547_ _04631_ memory\[35\]\[27\] _04617_ _04632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_191_4038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_191_4049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07098__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09478_ _03140_ _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07601__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08429_ _04011_ _01444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_210_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11123__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11440_ _05655_ _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_62_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_306_clk_i clknet_5_11__leaf_clk_i clknet_leaf_306_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_163_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10962__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11371_ _03311_ memory\[62\]\[1\] _05616_ _05618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13110_ memory\[20\]\[22\] memory\[21\]\[22\] _02368_ _02506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10322_ _05057_ _00211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14090_ _01129_ clknet_leaf_225_clk_i memory\[63\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12462__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13041_ memory\[22\]\[21\] memory\[23\]\[21\] _06751_ _02438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10253_ _05010_ memory\[46\]\[2\] _05006_ _05011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07048__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12697__A4 _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10184_ _04581_ memory\[45\]\[3\] _04969_ _04973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_167_3597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10952__I1 _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12529__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14992_ _02031_ clknet_leaf_62_clk_i memory\[38\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09263__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13943_ _00982_ clknet_leaf_130_clk_i memory\[8\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12854__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13874_ _00913_ clknet_leaf_61_clk_i memory\[39\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15613_ _00572_ clknet_leaf_333_clk_i memory\[58\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12825_ _06607_ _02224_ _02086_ _02225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_158_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10468__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15544_ _00503_ clknet_leaf_384_clk_i memory\[55\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12756_ memory\[16\]\[17\] memory\[17\]\[17\] memory\[18\]\[17\] memory\[19\]\[17\]
+ _06342_ _06485_ _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__12637__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07511__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11707_ _05689_ _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_7_Left_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15475_ _00434_ clknet_leaf_262_clk_i memory\[53\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12687_ _06610_ _02088_ _02089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14426_ _01465_ clknet_leaf_26_clk_i memory\[20\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09086__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11638_ memory\[24\]\[1\] memory\[25\]\[1\] memory\[26\]\[1\] memory\[27\]\[1\] _05778_
+ _05779_ _05853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13031__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14357_ _01396_ clknet_leaf_103_clk_i memory\[18\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11569_ _05784_ _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13308_ _02700_ net57 _02382_ _02701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08342__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14288_ _01327_ clknet_leaf_92_clk_i memory\[29\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_90_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13239_ _02371_ _02632_ _02373_ _02633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_412_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07800_ _03660_ _01166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08780_ _04202_ _01604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_127_Right_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07980__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09173__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07731_ _03184_ memory\[63\]\[19\] _03614_ _03624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09010__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11648__A2 _05855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11208__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07662_ _03587_ _01101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10112__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09401_ _04189_ memory\[34\]\[3\] _04538_ _04542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_172_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07593_ _03550_ _01069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09332_ _04505_ _01853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_66_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08517__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09263_ _04187_ memory\[32\]\[2\] _04466_ _04469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08214_ _03760_ memory\[17\]\[4\] _03893_ _03898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09194_ _04432_ _01788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12456__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08145_ _03861_ _01310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10782__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11584__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09348__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08252__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_84_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08076_ _03760_ memory\[15\]\[4\] _03819_ _03824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_292_clk_i clknet_5_15__leaf_clk_i clknet_leaf_292_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07027_ _03226_ _03117_ _03123_ _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_113_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08051__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10934__I1 _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08986__I _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12502__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08978_ _04317_ _01687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07929_ _03175_ memory\[19\]\[16\] _03722_ _03729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09001__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10022__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10940_ memory\[55\]\[23\] _03196_ _05385_ _05389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_230_clk_i clknet_5_26__leaf_clk_i clknet_leaf_230_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07563__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10871_ _05054_ memory\[54\]\[23\] _05348_ _05352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12610_ _06610_ _06810_ _06811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13261__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13590_ _05768_ _02973_ _02975_ _02977_ _02978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_66_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12541_ _06742_ _06743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_164_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_245_clk_i clknet_5_26__leaf_clk_i clknet_leaf_245_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_361_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08226__I _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15260_ _00219_ clknet_leaf_420_clk_i memory\[47\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12472_ _06610_ _06674_ _06675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_87_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11788__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14211_ _01250_ clknet_leaf_284_clk_i memory\[12\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11423_ _03363_ memory\[62\]\[26\] _05638_ _05645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15191_ _00150_ clknet_leaf_17_clk_i memory\[44\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12998__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11354_ _05608_ _00692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14142_ _01181_ clknet_leaf_285_clk_i memory\[7\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_169_3637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_89_Left_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10305_ _05045_ memory\[46\]\[19\] _05027_ _05046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_186_3951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14073_ _01112_ clknet_leaf_134_clk_i memory\[10\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11285_ _05571_ _00660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10236_ _04633_ memory\[45\]\[28\] _04991_ _05000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13024_ memory\[44\]\[21\] memory\[45\]\[21\] _02210_ _02421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11878__A2 _06088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10925__I1 _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13508__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09791__I1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10167_ _04963_ _00150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12827__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14975_ _02014_ clknet_leaf_421_clk_i memory\[38\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10098_ _04631_ memory\[43\]\[27\] _04919_ _04927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11028__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10689__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13926_ _00965_ clknet_leaf_212_clk_i memory\[8\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_98_Left_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13857_ _00896_ clknet_leaf_419_clk_i memory\[39\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10867__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12808_ _06446_ _02202_ _02204_ _02207_ _02208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__13252__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12686__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13788_ _00827_ clknet_leaf_371_clk_i memory\[16\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15527_ _00486_ clknet_leaf_289_clk_i memory\[55\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12739_ memory\[46\]\[17\] memory\[47\]\[17\] _06596_ _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09059__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15458_ _00417_ clknet_leaf_315_clk_i memory\[53\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07482__A2 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_61_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_106_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14409_ _01448_ clknet_leaf_189_clk_i memory\[20\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15389_ _00348_ clknet_leaf_347_clk_i memory\[51\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11566__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08072__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13307__A2 _02669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09950_ _04619_ memory\[41\]\[21\] _04847_ _04849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08901_ _04233_ memory\[26\]\[24\] _04272_ _04277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09881_ _04812_ _00015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13418__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08832_ _04237_ memory\[25\]\[26\] _04225_ _04238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09782__I1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07793__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07416__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08763_ _03137_ _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_139_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07714_ _03615_ _01125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13491__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08694_ _04152_ _01568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09631__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_140_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07645_ _03156_ memory\[10\]\[10\] _03578_ _03579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07170__A1 _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13153__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13243__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07576_ _03156_ memory\[0\]\[10\] _03541_ _03542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_101_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09298__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12277__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09315_ _04239_ memory\[32\]\[27\] _04488_ _04496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10852__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09246_ _04459_ _01813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_2_1_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_160_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09177_ _04237_ memory\[30\]\[26\] _04416_ _04423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08128_ _03812_ memory\[15\]\[29\] _03841_ _03851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09078__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10604__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09470__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08059_ _03813_ _01272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_147_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput46 net46 data_o[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_11070_ _05047_ memory\[57\]\[20\] _05457_ _05458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput57 net57 data_o[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09222__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08710__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput68 net68 data_o[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_11_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12601__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_308_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12740__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10021_ _04886_ _00081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07326__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output58_I net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14760_ _01799_ clknet_leaf_131_clk_i memory\[31\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11972_ memory\[44\]\[6\] memory\[45\]\[6\] _05749_ _06182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_153_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09541__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11332__I1 _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13711_ _03329_ memory\[9\]\[10\] _03086_ _03087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10923_ memory\[55\]\[15\] _03171_ _05374_ _05380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14691_ _01730_ clknet_leaf_358_clk_i memory\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10687__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_19_Right_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13642_ memory\[6\]\[31\] memory\[7\]\[31\] _05795_ _03029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_184_clk_i clknet_5_29__leaf_clk_i clknet_leaf_184_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13234__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10854_ _05037_ memory\[54\]\[15\] _05337_ _05343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12668__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07061__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11096__I0 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13573_ memory\[48\]\[30\] memory\[49\]\[30\] memory\[50\]\[30\] memory\[51\]\[30\]
+ _05725_ _05726_ _02961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10785_ _05306_ _00425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15312_ _00271_ clknet_leaf_158_clk_i memory\[48\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12524_ memory\[36\]\[14\] memory\[37\]\[14\] _06447_ _06726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15243_ _00202_ clknet_leaf_275_clk_i memory\[46\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_199_clk_i clknet_5_30__leaf_clk_i clknet_leaf_199_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12455_ _06450_ _06657_ _06177_ _06658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_140_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11311__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11548__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11406_ _03346_ memory\[62\]\[18\] _05627_ _05636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15174_ _00133_ clknet_leaf_32_clk_i memory\[44\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12386_ _06450_ _06589_ _06177_ _06590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XPHY_EDGE_ROW_28_Right_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14125_ _01164_ clknet_leaf_220_clk_i memory\[6\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12760__A3 _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11337_ _05599_ _00684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_122_clk_i clknet_5_23__leaf_clk_i clknet_leaf_122_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14056_ _01095_ clknet_leaf_215_clk_i memory\[10\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11268_ _05562_ _00652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12650__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13238__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13007_ _06851_ _02403_ _02404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11020__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12142__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10219_ _04968_ _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_11199_ _03344_ memory\[5\]\[17\] _05518_ _05526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_158_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07236__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09515__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_137_clk_i clknet_5_22__leaf_clk_i clknet_leaf_137_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11981__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_32_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14958_ _01997_ clknet_leaf_64_clk_i memory\[37\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_37_Right_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09451__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13909_ _00948_ clknet_leaf_113_clk_i memory\[11\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14889_ _01928_ clknet_leaf_47_clk_i memory\[35\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07430_ memory\[49\]\[7\] _03323_ _03455_ _03463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12028__A2 _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12659__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12097__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07361_ _03424_ _00963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09100_ _04382_ _01744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_21_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07292_ memory\[11\]\[8\] _03325_ _03379_ _03388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12825__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09031_ _04227_ memory\[28\]\[21\] _04344_ _04346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_257_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_46_Right_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09933_ _04602_ memory\[41\]\[13\] _04836_ _04840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08530__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09904__A1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09864_ _04803_ _00007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11711__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08815_ _04226_ _01615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_142_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09795_ memory\[3\]\[13\] _03165_ _04762_ _04766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12987__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11891__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_55_Right_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06985__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08746_ _04179_ _01593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13464__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13391__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_120_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08677_ memory\[23\]\[30\] _03371_ _04109_ _04143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07628_ _03132_ memory\[10\]\[2\] _03567_ _03570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11078__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07559_ _03132_ memory\[0\]\[2\] _03530_ _03533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11778__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_181_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10825__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10570_ _05180_ _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_106_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09691__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_64_Right_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_17_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09229_ _04450_ _01805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_118_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11131__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12240_ _05653_ _06446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_161_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09443__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12171_ _05699_ _06370_ _06377_ _06378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__11250__I0 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10970__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10753__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11122_ _05485_ _00583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_131_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12470__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11002__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13058__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_54_clk_i clknet_5_19__leaf_clk_i clknet_leaf_54_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11053_ _05031_ memory\[57\]\[12\] _05446_ _05449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06959__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12050__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_73_Right_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10004_ _04877_ _00073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14812_ _01851_ clknet_leaf_426_clk_i memory\[33\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15792_ _00751_ clknet_leaf_88_clk_i net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06895__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11305__I1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09271__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_69_clk_i clknet_5_16__leaf_clk_i clknet_leaf_69_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14743_ _01782_ clknet_leaf_86_clk_i memory\[30\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11955_ _06155_ _06158_ _06161_ _06164_ _06165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_28_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08182__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10906_ memory\[55\]\[7\] _03146_ _05363_ _05371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14674_ _01713_ clknet_leaf_83_clk_i memory\[28\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11886_ _06028_ _06096_ _05722_ _06097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13625_ memory\[60\]\[31\] memory\[61\]\[31\] _05702_ _03012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10837_ _05020_ memory\[54\]\[7\] _05326_ _05334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_82_Right_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_104_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13521__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13556_ _02375_ _02944_ _02945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_55_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10768_ _05297_ _00417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08615__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11864__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12507_ _03120_ _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13487_ _02494_ _02872_ _02874_ _02876_ _02877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_124_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10699_ _05018_ memory\[52\]\[6\] _05254_ _05261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15226_ _00185_ clknet_leaf_445_clk_i memory\[45\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12438_ _06640_ _06641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09434__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15157_ _00116_ clknet_leaf_10_clk_i memory\[43\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12369_ memory\[6\]\[12\] memory\[7\]\[12\] _06431_ _06573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07996__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14108_ _01147_ clknet_leaf_284_clk_i memory\[6\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08350__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13476__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15088_ _00047_ clknet_leaf_8_clk_i memory\[41\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_56_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_91_Right_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14039_ _01078_ clknet_leaf_54_clk_i memory\[0\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06930_ _03152_ _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_56_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07748__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input1_I address_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08600_ _03806_ memory\[22\]\[26\] _04095_ _04102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09580_ _04651_ _01955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13446__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09181__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08531_ _04065_ _01492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08173__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11216__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_6__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08462_ _03804_ memory\[20\]\[25\] _04023_ _04029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07413_ _03451_ _03452_ _03453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_08393_ _03992_ _01427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07344_ _03111_ memory\[8\]\[0\] _03415_ _03416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10807__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09673__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07275_ _03378_ _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_72_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09014_ _04210_ memory\[28\]\[13\] _04333_ _04337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12185__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11232__I0 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10790__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12280__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07987__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09356__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08260__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09916_ _04585_ memory\[41\]\[5\] _04825_ _04831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13685__A1 _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09847_ _04794_ _02079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11791__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09778_ memory\[3\]\[5\] _03140_ _04751_ _04757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08729_ _03798_ memory\[24\]\[22\] _04168_ _04171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11740_ memory\[6\]\[3\] memory\[7\]\[3\] _05706_ _05953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10030__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12660__A2 _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_83_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11671_ _05705_ _05884_ _05708_ _05885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13296__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13410_ memory\[44\]\[27\] memory\[45\]\[27\] _02210_ _02801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10622_ _05220_ _00348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08435__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14390_ _01429_ clknet_leaf_55_clk_i memory\[1\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09664__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13341_ _02732_ _02733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_172_3688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10553_ _05183_ _00316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_133_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13272_ _05772_ _02664_ _02195_ _02665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_162_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09416__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10484_ _05008_ memory\[4\]\[1\] _05145_ _05147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15011_ _02050_ clknet_leaf_339_clk_i memory\[3\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11796__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12223_ memory\[4\]\[10\] memory\[5\]\[10\] _06156_ _06429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07978__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12154_ _06149_ _06360_ _06361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_20_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11105_ _05476_ _00575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10205__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12479__A2 _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12085_ memory\[4\]\[8\] memory\[5\]\[8\] _06156_ _06293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13676__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_205_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11036_ _05014_ memory\[57\]\[4\] _05435_ _05440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_34_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13516__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13428__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12420__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15775_ _00734_ clknet_leaf_348_clk_i net65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12987_ memory\[60\]\[21\] memory\[61\]\[21\] _02164_ _02384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11036__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12100__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14726_ _01765_ clknet_leaf_132_clk_i memory\[30\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11938_ _06146_ _06147_ _05687_ _06148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08409__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07902__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14657_ _01696_ clknet_leaf_414_clk_i memory\[28\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10875__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11869_ memory\[54\]\[5\] memory\[55\]\[5\] _05684_ _06080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_25_Left_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_39_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13608_ _02995_ _02996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_28_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14588_ _01627_ clknet_leaf_390_clk_i memory\[26\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11837__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13539_ _05682_ _02927_ _02352_ _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_54_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07060_ _03245_ _00841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09407__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12167__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11214__I0 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15209_ _00168_ clknet_leaf_32_clk_i memory\[45\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_93_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07983__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07969__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_93_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08080__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_54_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_34_Left_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07962_ _03110_ _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_10_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13667__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_71_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09701_ _04577_ memory\[38\]\[1\] _04714_ _04716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06913_ net34 _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_71_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07893_ _03709_ _01210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08394__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09632_ _04679_ _01979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07424__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09563_ _04573_ memory\[36\]\[0\] _04642_ _04643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08146__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08514_ _04056_ _01484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09494_ _04574_ _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09894__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_407_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_43_Left_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08445_ _03787_ memory\[20\]\[17\] _04012_ _04020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_137_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_74_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08376_ _03983_ _01419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13198__A3 _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07327_ _03406_ _00947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_1_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08054__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_154_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07258_ _03366_ _00918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_30_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07189_ memory\[39\]\[5\] _03319_ _03309_ _03320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11905__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_52_Left_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09086__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13370__A3 _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11629__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08621__I1 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12005__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13658__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09814__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12330__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12910_ _02170_ _02307_ _02308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11764__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13890_ _00929_ clknet_leaf_303_clk_i memory\[11\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12881__A2 _02279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07334__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12841_ memory\[60\]\[19\] memory\[61\]\[19\] _02164_ _02240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_79_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_61_Left_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15560_ _00519_ clknet_leaf_232_clk_i memory\[56\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12772_ memory\[56\]\[18\] memory\[57\]\[18\] memory\[58\]\[18\] memory\[59\]\[18\]
+ _06827_ _02171_ _02172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_139_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14511_ _01550_ clknet_leaf_175_clk_i memory\[23\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_174_3728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11723_ memory\[60\]\[3\] memory\[61\]\[3\] _05656_ _05936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15491_ _00450_ clknet_leaf_335_clk_i memory\[54\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10695__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14442_ _01481_ clknet_leaf_192_clk_i memory\[21\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08165__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09637__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11654_ _05661_ _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_181_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12397__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10605_ _05210_ _00341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14373_ _01412_ clknet_leaf_338_clk_i memory\[1\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11585_ _05698_ _05730_ _05766_ _05800_ _05801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_107_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13324_ _02302_ _02708_ _02715_ _02716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_52_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10536_ _05060_ memory\[4\]\[26\] _05167_ _05174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_162_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Left_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13255_ _02647_ _02648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XPHY_EDGE_ROW_108_Right_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10467_ _05137_ _00276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07509__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12206_ memory\[60\]\[10\] memory\[61\]\[10\] _06273_ _06412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13186_ memory\[62\]\[24\] memory\[63\]\[24\] _02448_ _02580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10398_ _05058_ memory\[47\]\[25\] _05095_ _05101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12137_ _05783_ _06339_ _06341_ _06344_ _06345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA_clkbuf_leaf_356_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09724__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12068_ _05659_ _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12321__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11019_ _05430_ _00535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15827_ _00786_ clknet_leaf_121_clk_i memory\[9\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08128__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15758_ _00717_ clknet_leaf_221_clk_i memory\[62\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08679__I1 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14709_ _01748_ clknet_leaf_58_clk_i memory\[2\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15689_ _00648_ clknet_leaf_234_clk_i memory\[60\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08230_ _03906_ _01350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08161_ _03775_ memory\[29\]\[11\] _03868_ _03870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_95_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07112_ _03274_ _00864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08092_ _03832_ _01286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07043_ _03236_ _00833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12325__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12235__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11994__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08994_ _04326_ _01694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07945_ _03737_ _01234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08367__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07876_ _03197_ memory\[7\]\[23\] _03697_ _03701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10174__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09615_ _04627_ memory\[36\]\[25\] _04664_ _04670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_80_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09546_ _03208_ _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__06993__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09867__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_191_4039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09477_ _04584_ _01919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11404__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08428_ _03770_ memory\[20\]\[9\] _04001_ _04011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_50_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08359_ _03974_ _01411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_11__f_clk_i clknet_2_1_0_clk_i clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11370_ _05617_ _00699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10321_ _05056_ memory\[46\]\[24\] _05048_ _05057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13040_ _02436_ _02437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10252_ _03131_ _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12551__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10183_ _04972_ _00157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_167_3587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09544__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12969__I _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14991_ _02030_ clknet_leaf_43_clk_i memory\[38\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_128_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08358__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13066__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_128_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13942_ _00981_ clknet_leaf_130_clk_i memory\[8\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06967__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07030__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13873_ _00912_ clknet_leaf_62_clk_i memory\[39\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15612_ _00571_ clknet_leaf_331_clk_i memory\[58\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12824_ memory\[30\]\[18\] memory\[31\]\[18\] _02084_ _02224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15543_ _00502_ clknet_leaf_42_clk_i memory\[55\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12755_ _06480_ _02155_ _06482_ _02156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08530__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11706_ _05918_ _05919_ _05775_ _05920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15474_ _00433_ clknet_leaf_264_clk_i memory\[53\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12686_ memory\[24\]\[16\] memory\[25\]\[16\] memory\[26\]\[16\] memory\[27\]\[16\]
+ _06472_ _06611_ _02088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_126_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_413_clk_i clknet_5_2__leaf_clk_i clknet_leaf_413_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14425_ _01464_ clknet_leaf_98_clk_i memory\[20\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11417__I0 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11637_ _05772_ _05851_ _05775_ _05852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_65_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14356_ _01395_ clknet_leaf_104_clk_i memory\[18\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11568_ _03120_ _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08623__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12790__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13307_ _02654_ _02669_ _02684_ _02699_ _02700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_24_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10519_ _05043_ memory\[4\]\[18\] _05156_ _05165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10640__I1 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14287_ _01326_ clknet_leaf_184_clk_i memory\[29\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_428_clk_i clknet_5_1__leaf_clk_i clknet_leaf_428_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_64_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13414__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11499_ _05675_ _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_0_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09518__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07239__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13238_ memory\[22\]\[24\] memory\[23\]\[24\] _05754_ _02632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_90_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11984__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13169_ _02498_ _02563_ _02086_ _02564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_0_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13484__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_108_Left_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07730_ _03623_ _01133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_102_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10156__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07021__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07661_ _03181_ memory\[10\]\[18\] _03578_ _03587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09400_ _04541_ _01885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13704__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07592_ _03181_ memory\[0\]\[18\] _03541_ _03550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12153__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07702__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09331_ _04187_ memory\[33\]\[2\] _04502_ _04505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_66_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_87_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_103_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07324__I1 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11224__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09262_ _04468_ _01820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Left_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11408__I0 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08213_ _03897_ _01342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09193_ _04185_ memory\[31\]\[1\] _04430_ _04432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12456__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07088__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08144_ _03758_ memory\[29\]\[3\] _03857_ _03861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11584__A2 _05782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_27_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12781__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12055__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10631__I1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08075_ _03823_ _01278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07149__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07026_ _03116_ _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_101_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08588__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_126_Left_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09364__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08977_ _04241_ memory\[27\]\[28\] _04308_ _04317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11693__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07928_ _03728_ _01226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10147__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07859_ _03172_ memory\[7\]\[15\] _03686_ _03692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13614__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_123_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10870_ _05351_ _00465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08708__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09529_ _04619_ memory\[35\]\[21\] _04617_ _04620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07315__I1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12540_ memory\[28\]\[14\] memory\[29\]\[14\] _06604_ _06742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_304_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12471_ memory\[24\]\[13\] memory\[25\]\[13\] memory\[26\]\[13\] memory\[27\]\[13\]
+ _06472_ _06611_ _06674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_19_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13644__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14210_ _01249_ clknet_leaf_282_clk_i memory\[12\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_193_Right_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11422_ _05644_ _00724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_191_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08443__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15190_ _00149_ clknet_leaf_16_clk_i memory\[44\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14141_ _01180_ clknet_leaf_286_clk_i memory\[7\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11353_ memory\[61\]\[25\] _03202_ _05602_ _05608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_169_3627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07059__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10304_ _03183_ _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_14072_ _01111_ clknet_leaf_134_clk_i memory\[10\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11284_ _03361_ memory\[60\]\[25\] _05565_ _05571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_186_3952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08579__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13023_ _02337_ _02415_ _02417_ _02419_ _02420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10235_ _04999_ _00182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10166_ _04631_ memory\[44\]\[27\] _04955_ _04963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10213__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14974_ _02013_ clknet_leaf_419_clk_i memory\[38\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10097_ _04926_ _00117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13925_ _00964_ clknet_leaf_298_clk_i memory\[8\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13856_ _00895_ clknet_leaf_418_clk_i memory\[39\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12135__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12807_ _06453_ _02206_ _02207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_130_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13787_ _00826_ clknet_leaf_394_clk_i memory\[14\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08503__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_352_clk_i clknet_5_8__leaf_clk_i clknet_leaf_352_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10999_ _05045_ memory\[56\]\[19\] _05410_ _05420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12686__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11044__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12738_ _02138_ _02139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15526_ _00485_ clknet_leaf_288_clk_i memory\[55\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_44_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_44_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15457_ _00416_ clknet_leaf_330_clk_i memory\[53\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10883__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12669_ _06453_ _06868_ _06869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_170_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14408_ _01447_ clknet_leaf_182_clk_i memory\[20\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09449__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_160_Right_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15388_ _00347_ clknet_leaf_346_clk_i memory\[51\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13479__B _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_367_clk_i clknet_5_9__leaf_clk_i clknet_leaf_367_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14339_ _01378_ clknet_leaf_342_clk_i memory\[18\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13307__A3 _02684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08900_ _04276_ _01650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09880_ _04616_ memory\[40\]\[20\] _04811_ _04812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10377__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08831_ _03205_ _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_08762_ _04190_ _01598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_253_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_305_clk_i clknet_5_11__leaf_clk_i clknet_leaf_305_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07713_ _03156_ memory\[63\]\[10\] _03614_ _03615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09912__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08693_ _03762_ memory\[24\]\[5\] _04146_ _04152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_105_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13434__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07644_ _03566_ _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08528__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07432__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_101_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07575_ _03529_ _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_101_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09314_ _04495_ _01845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07231__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09245_ _04237_ memory\[31\]\[26\] _04452_ _04459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09176_ _04422_ _01780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08127_ _03850_ _01303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_4_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08058_ _03812_ memory\[12\]\[29\] _03794_ _03813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12506__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput47 net47 data_o[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_07009_ _03212_ memory\[14\]\[28\] _03188_ _03213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13609__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput58 net58 data_o[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12513__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput69 net69 data_o[7] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09094__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12601__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07607__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10020_ _04621_ memory\[42\]\[22\] _04883_ _04886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11637__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11129__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08981__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_76_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09822__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10968__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11971_ _05732_ _06175_ _06178_ _06180_ _06181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08733__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__I1 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13710_ _03074_ _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11493__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10922_ _05379_ _00489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14690_ _01729_ clknet_leaf_360_clk_i memory\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10540__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13641_ _03027_ _03028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_156_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10853_ _05342_ _00457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12668__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_184_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13572_ _05719_ _02959_ _05739_ _02960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_82_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10784_ _05035_ memory\[53\]\[14\] _05301_ _05306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_742 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15311_ _00270_ clknet_leaf_256_clk_i memory\[48\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12993__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12523_ _06428_ _06712_ _06724_ _06725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_13_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09269__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15242_ _00201_ clknet_leaf_275_clk_i memory\[46\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08173__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06980__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12454_ memory\[38\]\[13\] memory\[39\]\[13\] _06039_ _06657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11405_ _05635_ _00716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15173_ _00132_ clknet_leaf_430_clk_i memory\[44\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12385_ memory\[38\]\[12\] memory\[39\]\[12\] _06039_ _06589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14124_ _01163_ clknet_leaf_220_clk_i memory\[6\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11336_ memory\[61\]\[17\] _03177_ _05591_ _05599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08901__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12760__A4 _02160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14055_ _01094_ clknet_leaf_212_clk_i memory\[10\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11267_ _03344_ memory\[60\]\[17\] _05554_ _05562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13006_ memory\[0\]\[21\] memory\[1\]\[21\] memory\[2\]\[21\] memory\[3\]\[21\] _06709_
+ _06779_ _02403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_24_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07517__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10218_ _04990_ _00174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11198_ _05525_ _00619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11720__A2 _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12222__I _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10149_ _04614_ memory\[44\]\[19\] _04944_ _04954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09732__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12356__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_85_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14957_ _01996_ clknet_leaf_49_clk_i memory\[37\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13254__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13908_ _00947_ clknet_leaf_129_clk_i memory\[11\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08348__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14888_ _01927_ clknet_leaf_46_clk_i memory\[35\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09531__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13839_ _00878_ clknet_leaf_197_clk_i memory\[13\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12659__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07360_ _03150_ memory\[8\]\[8\] _03415_ _03424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15509_ _00468_ clknet_leaf_155_clk_i memory\[54\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07291_ _03387_ _00930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07986__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09030_ _04345_ _01711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09179__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06890__I net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13528__A3 _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10118__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10598__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_170_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_106_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09932_ _04839_ _00039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12333__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09904__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09863_ _04600_ memory\[40\]\[12\] _04800_ _04803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08963__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_244_clk_i clknet_5_26__leaf_clk_i clknet_leaf_244_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08814_ _04224_ memory\[25\]\[20\] _04225_ _04226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_142_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09794_ _04765_ _02055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_77_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08745_ _03814_ memory\[24\]\[30\] _04145_ _04179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10788__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08258__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08676_ _04142_ _01560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_259_clk_i clknet_5_13__leaf_clk_i clknet_leaf_259_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_120_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08340__A1 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07627_ _03569_ _01084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08057__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07558_ _03532_ _01052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_157_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_180_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07489_ _03495_ _01020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09228_ _04220_ memory\[31\]\[18\] _04441_ _04450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_185_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12727__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09159_ _04413_ _01772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10028__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10589__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_135_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12170_ _06024_ _06372_ _06374_ _06376_ _06377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_102_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11121_ _03334_ memory\[58\]\[12\] _05482_ _05485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_131_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output70_I net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12586__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11052_ _05448_ _00550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08954__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10003_ _04604_ memory\[42\]\[14\] _04872_ _04877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10761__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14811_ _01850_ clknet_leaf_0_clk_i memory\[32\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12977__I _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15791_ _00750_ clknet_leaf_253_clk_i net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_98_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08706__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_149_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07509__I1 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06975__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14742_ _01781_ clknet_leaf_88_clk_i memory\[30\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11954_ _06162_ _06163_ _06164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_118_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10513__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07072__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10905_ _05370_ _00481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14673_ _01712_ clknet_leaf_91_clk_i memory\[28\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11885_ memory\[14\]\[5\] memory\[15\]\[5\] _05720_ _06096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13624_ _03011_ _00761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_184_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10836_ _05333_ _00449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12926__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09131__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13555_ memory\[16\]\[29\] memory\[17\]\[29\] memory\[18\]\[29\] memory\[19\]\[29\]
+ _05761_ _02376_ _02944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_66_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_201_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10767_ _05018_ memory\[53\]\[6\] _05290_ _05297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11322__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12506_ _06159_ _06706_ _06707_ _06708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13486_ _02501_ _02875_ _02876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_42_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10698_ _05260_ _00384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12718__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15225_ _00184_ clknet_leaf_23_clk_i memory\[45\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12437_ memory\[4\]\[13\] memory\[5\]\[13\] _06156_ _06640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_152_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13391__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_23_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15156_ _00115_ clknet_leaf_10_clk_i memory\[43\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12368_ _06571_ _06572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08631__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13249__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_39_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14107_ _01146_ clknet_leaf_389_clk_i memory\[63\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_39_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11319_ memory\[61\]\[9\] _03152_ _05580_ _05590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15087_ _00046_ clknet_leaf_19_clk_i memory\[41\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12299_ memory\[48\]\[11\] memory\[49\]\[11\] memory\[50\]\[11\] memory\[51\]\[11\]
+ _06010_ _06150_ _06504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08430__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14038_ _01077_ clknet_leaf_55_clk_i memory\[0\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_56_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11992__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12329__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_171_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08530_ _03804_ memory\[21\]\[25\] _04059_ _04065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11457__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06885__I net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08078__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08461_ _04028_ _01459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07412_ _03226_ _03117_ _03265_ _03452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_175_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08392_ _03802_ memory\[1\]\[24\] _03987_ _03992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07710__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12957__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07343_ _03414_ _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_85_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11232__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07684__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07274_ _03377_ _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09013_ _04336_ _01703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09637__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_76_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_76_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_403_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10991__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07157__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09436__I _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13134__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_183_clk_i clknet_5_29__leaf_clk_i clknet_leaf_183_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09915_ _04830_ _00031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13685__A2 _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12732__I1 memory\[39\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09846_ _04583_ memory\[40\]\[4\] _04789_ _04794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10743__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11791__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09777_ _04756_ _02047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06989_ _03197_ memory\[14\]\[23\] _03188_ _03198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_150_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_198_clk_i clknet_5_31__leaf_clk_i clknet_leaf_198_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08728_ _04170_ _01584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08659_ memory\[23\]\[21\] _03353_ _04132_ _04134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_159_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_121_clk_i clknet_5_23__leaf_clk_i clknet_leaf_121_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11670_ memory\[6\]\[2\] memory\[7\]\[2\] _05706_ _05884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08716__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09113__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13296__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10621_ memory\[51\]\[1\] _03128_ _05218_ _05220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11142__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_12_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13340_ memory\[36\]\[26\] memory\[37\]\[26\] _02338_ _02732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_172_3678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10552_ _05008_ memory\[50\]\[1\] _05181_ _05183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_172_3689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_136_clk_i clknet_5_22__leaf_clk_i clknet_leaf_136_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13748__I0 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13271_ memory\[14\]\[25\] memory\[15\]\[25\] _02193_ _02664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10981__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10483_ _05146_ _00283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15010_ _02049_ clknet_leaf_339_clk_i memory\[3\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12222_ _03114_ _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09547__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_75_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12153_ memory\[48\]\[9\] memory\[49\]\[9\] memory\[50\]\[9\] memory\[51\]\[9\] _06010_
+ _06150_ _06360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_102_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07067__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11104_ _03317_ memory\[58\]\[4\] _05471_ _05476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12084_ _05651_ _06283_ _06291_ _06292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_21_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08927__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11035_ _05439_ _00542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11687__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09282__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11317__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12986_ _02383_ _00751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15774_ _00733_ clknet_leaf_348_clk_i net62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09352__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14725_ _01764_ clknet_leaf_410_clk_i memory\[30\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_24_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11937_ memory\[54\]\[6\] memory\[55\]\[6\] _05684_ _06147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11116__I _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14656_ _01695_ clknet_leaf_413_clk_i memory\[28\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11868_ _06078_ _06079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07530__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11560__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10819_ _05070_ memory\[53\]\[31\] _05289_ _05324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13607_ memory\[28\]\[30\] memory\[29\]\[30\] _02495_ _02995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_352_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11799_ memory\[48\]\[4\] memory\[49\]\[4\] memory\[50\]\[4\] memory\[51\]\[4\] _06010_
+ _05694_ _06011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_14587_ _01626_ clknet_leaf_4_clk_i memory\[25\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_54_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07666__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13538_ memory\[46\]\[29\] memory\[47\]\[29\] _02487_ _02927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13469_ _02341_ _02858_ _05708_ _02859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_152_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09457__S _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15208_ _00167_ clknet_leaf_32_clk_i memory\[45\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_93_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08091__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15139_ _00098_ clknet_leaf_433_clk_i memory\[43\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13116__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07961_ _03745_ _01242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09700_ _04715_ _02011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06912_ _03139_ _00799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11678__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07892_ _03221_ memory\[7\]\[31\] _03674_ _03709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09631_ _04573_ memory\[37\]\[0\] _04678_ _04679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09562_ _04641_ _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10131__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09343__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08513_ _03787_ memory\[21\]\[17\] _04048_ _04056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09920__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09493_ _03155_ _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11150__I0 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08444_ _04019_ _01451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08536__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_4092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08375_ _03785_ memory\[1\]\[16\] _03976_ _03983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_163_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_53_clk_i clknet_5_19__leaf_clk_i clknet_leaf_53_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_154_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07326_ memory\[11\]\[24\] _03359_ _03401_ _03406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07657__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11602__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_115_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07257_ memory\[39\]\[27\] _03365_ _03351_ _03366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_30_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_30_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_68_clk_i clknet_5_16__leaf_clk_i clknet_leaf_68_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07188_ _03140_ _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08082__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10964__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08909__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10716__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07615__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12330__A2 _06534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11764__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09829_ _04783_ _02072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12840_ _02239_ _00749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09830__S _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12771_ _03116_ _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_55_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10976__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14510_ _01549_ clknet_leaf_174_clk_i memory\[23\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11722_ _05935_ _00733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_174_3718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15490_ _00449_ clknet_leaf_337_clk_i memory\[54\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07896__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_174_3729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07350__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14441_ _01480_ clknet_leaf_189_clk_i memory\[21\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11653_ _05866_ _05867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10775__I _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10604_ _05060_ memory\[50\]\[26\] _05203_ _05210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14372_ _01411_ clknet_leaf_281_clk_i memory\[1\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11584_ _05767_ _05782_ _05799_ _05800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_25_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13323_ _05715_ _02710_ _02712_ _02714_ _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10535_ _05173_ _00308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09277__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13254_ memory\[52\]\[25\] memory\[53\]\[25\] _06832_ _02647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10466_ _05058_ memory\[48\]\[25\] _05131_ _05137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07025__A1 _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12205_ _03450_ _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_32_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13185_ _02578_ _02579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_36_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10397_ _05100_ _00243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12136_ _05794_ _06343_ _06344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07820__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10015__I _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12067_ _06274_ _06275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12431__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07525__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09573__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11018_ _05064_ memory\[56\]\[28\] _05421_ _05430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_189_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15826_ _00785_ clknet_leaf_122_clk_i memory\[9\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12704__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15757_ _00716_ clknet_leaf_224_clk_i memory\[62\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12969_ _05747_ _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__13262__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14708_ _01747_ clknet_leaf_57_clk_i memory\[2\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_16_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08356__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11832__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15688_ _00647_ clknet_leaf_236_clk_i memory\[60\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12386__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07260__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14639_ _01678_ clknet_leaf_125_clk_i memory\[27\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08160_ _03869_ _01317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_95_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07111_ _03141_ memory\[13\]\[5\] _03268_ _03274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08091_ _03775_ memory\[15\]\[11\] _03830_ _03832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13337__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09187__S _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07042_ _03144_ memory\[16\]\[6\] _03229_ _03236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08091__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11199__I0 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10126__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08064__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_110_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11994__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08993_ _04189_ memory\[28\]\[3\] _04322_ _04326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07944_ _03197_ memory\[19\]\[23\] _03733_ _03737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07875_ _03700_ _01201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11371__I0 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_3_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09614_ _04669_ _01971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_23_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07234__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13680__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09545_ _04630_ _01941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_151_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11123__I0 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_174_Right_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07878__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09476_ _04583_ memory\[35\]\[4\] _04575_ _04584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11823__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08266__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08427_ _04010_ _01443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13576__A1 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08358_ _03768_ memory\[1\]\[8\] _03965_ _03974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_248_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07309_ memory\[11\]\[16\] _03342_ _03390_ _03397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12516__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08289_ _03937_ _01378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13328__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09097__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10320_ _03199_ _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_14_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08055__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10251_ _05009_ _00188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10036__S _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10182_ _04579_ memory\[45\]\[2\] _04969_ _04972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_300_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_167_3599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13347__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14990_ _02029_ clknet_leaf_43_clk_i memory\[38\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_31_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12934__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13941_ _00980_ clknet_leaf_129_clk_i memory\[8\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13872_ _00911_ clknet_leaf_61_clk_i memory\[39\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_9_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09307__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15611_ _00570_ clknet_leaf_376_clk_i memory\[57\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12823_ _02222_ _02223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_119_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11114__I0 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13082__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_141_Right_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06983__I net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15542_ _00501_ clknet_leaf_42_clk_i memory\[55\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12754_ memory\[22\]\[17\] memory\[23\]\[17\] _06751_ _02155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07080__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11705_ memory\[30\]\[2\] memory\[31\]\[2\] _05773_ _05919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12685_ _06607_ _02085_ _02086_ _02087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_126_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15473_ _00432_ clknet_leaf_261_clk_i memory\[53\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13567__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14424_ _01463_ clknet_leaf_92_clk_i memory\[20\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11636_ memory\[30\]\[1\] memory\[31\]\[1\] _05773_ _05851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_65_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14355_ _01394_ clknet_leaf_101_clk_i memory\[18\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11567_ _05747_ _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11330__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13306_ _02358_ _02691_ _02698_ _02699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10518_ _05164_ _00300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14286_ _01325_ clknet_leaf_183_clk_i memory\[29\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08703__I _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11498_ _05700_ _05704_ _05709_ _05713_ _05714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_150_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13414__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08046__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13237_ _02630_ _02631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_90_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12225__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10449_ _05041_ memory\[48\]\[17\] _05120_ _05128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13168_ memory\[30\]\[23\] memory\[31\]\[23\] _02084_ _02563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12119_ memory\[40\]\[8\] memory\[41\]\[8\] memory\[42\]\[8\] memory\[43\]\[8\] _06186_
+ _06326_ _06327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
X_13099_ _05655_ _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_97_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09534__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07660_ _03586_ _01100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09470__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_197_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12058__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15809_ _00768_ clknet_leaf_301_clk_i memory\[9\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07591_ _03549_ _01068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09330_ _04504_ _01852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07989__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11505__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12153__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08086__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09261_ _04185_ memory\[32\]\[1\] _04466_ _04468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13005__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13558__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08212_ _03758_ memory\[17\]\[3\] _03893_ _03897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09192_ _04431_ _01787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08814__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12844__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08143_ _03860_ _01309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12230__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11664__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11240__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10092__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08985__A1 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08074_ _03758_ memory\[15\]\[3\] _03819_ _03823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08037__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07025_ _03112_ _03224_ _03225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_60_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_149_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09645__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07260__I1 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08976_ _04316_ _01686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input32_I data_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07165__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07927_ _03172_ memory\[19\]\[15\] _03722_ _03728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_162_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07858_ _03691_ _01193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12049__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07789_ _03169_ memory\[6\]\[14\] _03650_ _03655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11415__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09528_ _03190_ _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_78_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13261__A3 _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09459_ _04247_ memory\[34\]\[31\] _04537_ _04572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13549__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12470_ _06607_ _06672_ _06195_ _06673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_136_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_35_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_399_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11421_ _03361_ memory\[62\]\[25\] _05638_ _05644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13644__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08276__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12221__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11150__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14140_ _01179_ clknet_leaf_284_clk_i memory\[7\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11352_ _05607_ _00691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10303_ _05044_ _00205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14071_ _01110_ clknet_leaf_135_clk_i memory\[10\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11283_ _05570_ _00659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_186_3953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13022_ _02344_ _02418_ _02419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_162_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10234_ _04631_ memory\[45\]\[27\] _04991_ _04999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10165_ _04962_ _00149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07251__I1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14973_ _02012_ clknet_leaf_427_clk_i memory\[38\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10096_ _04629_ memory\[43\]\[26\] _04919_ _04926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08200__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13924_ _00963_ clknet_leaf_299_clk_i memory\[8\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09290__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13855_ _00894_ clknet_leaf_419_clk_i memory\[39\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12135__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12806_ memory\[32\]\[18\] memory\[33\]\[18\] memory\[34\]\[18\] memory\[35\]\[18\]
+ _02205_ _06454_ _02206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_97_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13786_ _00825_ clknet_leaf_386_clk_i memory\[14\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10998_ _05419_ _00525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15525_ _00484_ clknet_leaf_312_clk_i memory\[55\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12737_ memory\[44\]\[17\] memory\[45\]\[17\] _06319_ _02138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_44_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15456_ _00415_ clknet_leaf_330_clk_i memory\[53\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12668_ memory\[32\]\[16\] memory\[33\]\[16\] memory\[34\]\[16\] memory\[35\]\[16\]
+ _06314_ _06454_ _06868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_154_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_61_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14407_ _01446_ clknet_leaf_190_clk_i memory\[20\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11619_ memory\[36\]\[1\] memory\[37\]\[1\] _05733_ _05834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12212__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15387_ _00346_ clknet_leaf_378_clk_i memory\[50\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12599_ memory\[46\]\[15\] memory\[47\]\[15\] _06596_ _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_167_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14338_ _01377_ clknet_leaf_341_clk_i memory\[18\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13399__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_40_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07490__I1 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14269_ _01308_ clknet_leaf_390_clk_i memory\[29\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08830_ _04236_ _01620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07242__I1 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10404__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09519__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08761_ _04189_ memory\[25\]\[3\] _04183_ _04190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13715__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07712_ _03602_ _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_100_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08692_ _04151_ _01567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_68_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07713__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07643_ _03577_ _01092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_140_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07574_ _03540_ _01060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13243__A3 _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09313_ _04237_ memory\[32\]\[26\] _04488_ _04495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12451__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09244_ _04458_ _01812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_7_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08258__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09175_ _04235_ memory\[30\]\[25\] _04416_ _04422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12066__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10065__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08126_ _03810_ memory\[15\]\[28\] _03841_ _03850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Right_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08057_ _03214_ _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07008_ _03211_ _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09375__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput48 net48 data_o[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput59 net59 data_o[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_164_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_412_clk_i clknet_5_2__leaf_clk_i clknet_leaf_412_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_181_3861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08959_ _04307_ _01678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13625__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11970_ _05741_ _06179_ _06180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_93_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_5_26__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10921_ memory\[55\]\[14\] _03168_ _05374_ _05379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11493__A2 _05707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_427_clk_i clknet_5_2__leaf_clk_i clknet_leaf_427_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_169_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13314__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13640_ memory\[4\]\[31\] memory\[5\]\[31\] _05789_ _03027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10852_ _05035_ memory\[54\]\[14\] _05337_ _05342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12442__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13571_ memory\[54\]\[30\] memory\[55\]\[30\] _05720_ _02959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10783_ _05305_ _00424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_186_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15310_ _00269_ clknet_leaf_256_clk_i memory\[48\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12522_ _06713_ _06716_ _06719_ _06723_ _06724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_137_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08454__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11879__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15241_ _00200_ clknet_leaf_277_clk_i memory\[46\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12453_ _06655_ _06656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10056__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11404_ _03344_ memory\[62\]\[17\] _05627_ _05635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_145_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09997__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15172_ _00131_ clknet_leaf_399_clk_i memory\[44\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12384_ _06587_ _06588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_34_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14123_ _01162_ clknet_leaf_221_clk_i memory\[6\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07621__A1 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11335_ _05598_ _00683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07472__I1 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09749__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14054_ _01093_ clknet_leaf_216_clk_i memory\[10\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11266_ _05561_ _00651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13005_ _06848_ _02401_ _06707_ _02402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10217_ _04614_ memory\[45\]\[19\] _04980_ _04990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10224__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11197_ _03342_ memory\[5\]\[16\] _05518_ _05525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11720__A3 _05913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10148_ _04953_ _00141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12356__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10079_ _04612_ memory\[43\]\[18\] _04908_ _04917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_85_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14956_ _01995_ clknet_leaf_48_clk_i memory\[37\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08629__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_145_Left_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13907_ _00946_ clknet_leaf_120_clk_i memory\[11\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14887_ _01926_ clknet_leaf_49_clk_i memory\[35\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11055__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13838_ _00877_ clknet_leaf_196_clk_i memory\[13\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_63_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10894__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08488__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13769_ _00808_ clknet_leaf_217_clk_i memory\[14\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_21_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15508_ _00467_ clknet_leaf_155_clk_i memory\[54\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07290_ memory\[11\]\[7\] _03323_ _03379_ _03387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12394__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11789__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15439_ _00398_ clknet_leaf_274_clk_i memory\[52\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_154_Left_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09988__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12292__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12614__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09195__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07708__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09931_ _04600_ memory\[41\]\[12\] _04836_ _04839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_146_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08412__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09862_ _04802_ _00006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_347_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08813_ _04182_ _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_142_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_142_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09793_ memory\[3\]\[12\] _03162_ _04762_ _04765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_163_Left_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13445__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08744_ _04178_ _01592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07443__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12569__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09912__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08675_ memory\[23\]\[29\] _03369_ _04132_ _04142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_120_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07626_ _03129_ memory\[10\]\[1\] _03567_ _03569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07557_ _03129_ memory\[0\]\[1\] _03530_ _03532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_187_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07488_ memory\[59\]\[1\] _03311_ _03493_ _03495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08274__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07151__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_172_Left_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09227_ _04449_ _01804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10309__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10038__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09158_ _04218_ memory\[30\]\[17\] _04405_ _04413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12727__A2 _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08109_ _03818_ _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_133_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09089_ _04376_ _01739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12524__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11120_ _05484_ _00582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_183_3901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12035__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11051_ _05029_ memory\[57\]\[11\] _05446_ _05448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12586__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10044__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_351_clk_i clknet_5_8__leaf_clk_i clknet_leaf_351_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output63_I net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_181_Left_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10002_ _04876_ _00072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13355__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14810_ _01849_ clknet_leaf_5_clk_i memory\[32\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08449__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15790_ _00749_ clknet_leaf_253_clk_i net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_157_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_366_clk_i clknet_5_9__leaf_clk_i clknet_leaf_366_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14741_ _01780_ clknet_leaf_87_clk_i memory\[30\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11953_ memory\[0\]\[6\] memory\[1\]\[6\] memory\[2\]\[6\] memory\[3\]\[6\] _06020_
+ _06090_ _06163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_192_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_169_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_71_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10904_ memory\[55\]\[6\] _03143_ _05363_ _05370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14672_ _01711_ clknet_leaf_91_clk_i memory\[28\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07390__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11884_ _06094_ _06095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_169_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13623_ _03010_ net63 _03122_ _03011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10835_ _05018_ memory\[54\]\[6\] _05326_ _05333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06893__A2 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_190_Left_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06991__I net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13554_ _02371_ _02942_ _02373_ _02943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08184__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10766_ _05296_ _00416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12505_ _05686_ _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_125_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08890__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13485_ memory\[24\]\[28\] memory\[25\]\[28\] memory\[26\]\[28\] memory\[27\]\[28\]
+ _02363_ _02502_ _02875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10697_ _05016_ memory\[52\]\[5\] _05254_ _05260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12718__A2 _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_304_clk_i clknet_5_11__leaf_clk_i clknet_leaf_304_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15224_ _00183_ clknet_leaf_23_clk_i memory\[45\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_296_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12436_ _06411_ _06631_ _06638_ _06639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_120_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15155_ _00114_ clknet_leaf_11_clk_i memory\[43\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07445__I1 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12367_ memory\[4\]\[12\] memory\[5\]\[12\] _06156_ _06571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07528__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14106_ _01145_ clknet_leaf_387_clk_i memory\[63\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_39_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11318_ _05589_ _00675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15086_ _00045_ clknet_leaf_20_clk_i memory\[41\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12298_ _06146_ _06502_ _06287_ _06503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_319_clk_i clknet_5_11__leaf_clk_i clknet_leaf_319_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14037_ _01076_ clknet_leaf_56_clk_i memory\[0\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11249_ _05552_ _00643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10201__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09743__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06956__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12329__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07263__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12654__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14939_ _01978_ clknet_leaf_444_clk_i memory\[36\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08460_ _03802_ memory\[20\]\[24\] _04023_ _04028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08158__I _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07381__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07411_ _03112_ _03450_ _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_174_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08391_ _03991_ _01426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10268__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07342_ _03115_ net73 _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_163_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12957__A2 _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07273_ _03115_ _03376_ _03377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_TAPCELL_ROW_14_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09012_ _04208_ memory\[28\]\[12\] _04333_ _04336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_143_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_76_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_76_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09914_ _04583_ memory\[41\]\[4\] _04825_ _04830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09845_ _04793_ _02078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10799__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13175__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09776_ memory\[3\]\[4\] _03137_ _04751_ _04756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06988_ _03196_ _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08727_ _03796_ memory\[24\]\[21\] _04168_ _04170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08658_ _04133_ _01551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_159_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07609_ _03206_ memory\[0\]\[26\] _03552_ _03559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08589_ _04096_ _01519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_176_3760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_176_3771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11423__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10259__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10620_ _05219_ _00347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07124__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_12_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10551_ _05182_ _00315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08872__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_172_3679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09828__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13270_ _02662_ _02663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10482_ _05004_ memory\[4\]\[0\] _05145_ _05146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_18_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12221_ _06411_ _06418_ _06426_ _06427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__12254__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12420__I1 net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07348__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12152_ _06146_ _06358_ _06287_ _06359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_124_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_290_clk_i clknet_5_15__leaf_clk_i clknet_leaf_290_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11103_ _05475_ _00574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12083_ _06142_ _06285_ _06288_ _06290_ _06291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_60_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09563__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11034_ _05012_ memory\[57\]\[3\] _05435_ _05439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12884__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_188_Right_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_5_2__f_clk_i clknet_2_0_0_clk_i clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_51_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15773_ _00732_ clknet_leaf_342_clk_i net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12985_ _02381_ net52 _02382_ _02383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10498__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14724_ _01763_ clknet_leaf_405_clk_i memory\[30\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10301__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11936_ _05681_ _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08907__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14655_ _01694_ clknet_leaf_354_clk_i memory\[28\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11867_ memory\[52\]\[5\] memory\[53\]\[5\] _05678_ _06078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12429__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_156_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13606_ _03304_ _02986_ _02993_ _02994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_156_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10818_ _05323_ _00441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13061__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14586_ _01625_ clknet_leaf_3_clk_i memory\[25\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07115__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11798_ _05691_ _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_171_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_27_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13537_ _02925_ _02926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_243_clk_i clknet_5_26__leaf_clk_i clknet_leaf_243_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_171_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08863__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10749_ _05068_ memory\[52\]\[30\] _05253_ _05287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09738__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13468_ memory\[38\]\[28\] memory\[39\]\[28\] _05662_ _02858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15207_ _00166_ clknet_leaf_31_clk_i memory\[45\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07418__I1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12419_ _06570_ _06586_ _06602_ _06622_ _06623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__12164__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13399_ memory\[8\]\[27\] memory\[9\]\[27\] memory\[10\]\[27\] memory\[11\]\[27\]
+ _02473_ _05779_ _02790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_26_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09537__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10422__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_258_clk_i clknet_5_13__leaf_clk_i clknet_leaf_258_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15138_ _00097_ clknet_leaf_442_clk_i memory\[43\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15069_ _00028_ clknet_leaf_434_clk_i memory\[41\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07960_ _03221_ memory\[19\]\[31\] _03710_ _03745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09473__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06911_ _03138_ memory\[14\]\[4\] _03126_ _03139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_71_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07891_ _03708_ _01209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_155_Right_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09630_ _04677_ _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08089__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09561_ _03305_ _03750_ _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__13723__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08512_ _04055_ _01483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08817__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09492_ _04594_ _01924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07354__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07721__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08443_ _03785_ memory\[20\]\[16\] _04012_ _04019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_193_4093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_137_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08374_ _03982_ _01418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07325_ _03405_ _00946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_154_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07256_ _03208_ _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_115_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08552__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08606__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07187_ _03318_ _00895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_182_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09383__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09031__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12866__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_122_Right_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09828_ memory\[3\]\[29\] _03214_ _04773_ _04783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_244_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09759_ _04635_ memory\[38\]\[29\] _04736_ _04746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12770_ _05667_ _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__13291__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08727__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11721_ _05934_ net62 _05802_ _05935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_174_3719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14440_ _01479_ clknet_leaf_182_clk_i memory\[21\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11652_ memory\[60\]\[2\] memory\[61\]\[2\] _05656_ _05866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_182_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10603_ _05209_ _00340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14371_ _01410_ clknet_leaf_339_clk_i memory\[1\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11583_ _05783_ _05787_ _05793_ _05798_ _05799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_37_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13322_ _05724_ _02713_ _02714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08462__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10534_ _05058_ memory\[4\]\[25\] _05167_ _05173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07273__A2 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_49_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13253_ _02163_ _02641_ _02643_ _02645_ _02646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10465_ _05136_ _00275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_20_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12204_ _06410_ _00740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10404__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07025__A2 _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13184_ memory\[60\]\[24\] memory\[61\]\[24\] _02164_ _02578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10396_ _05056_ memory\[47\]\[24\] _05095_ _05100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12135_ memory\[16\]\[8\] memory\[17\]\[8\] memory\[18\]\[8\] memory\[19\]\[8\] _06342_
+ _05796_ _06343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_20_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_53_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07806__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09022__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11836__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12066_ memory\[60\]\[8\] memory\[61\]\[8\] _06273_ _06274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11328__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12511__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11017_ _05429_ _00534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10232__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15825_ _00784_ clknet_leaf_128_clk_i memory\[9\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15756_ _00715_ clknet_leaf_223_clk_i memory\[62\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12704__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12968_ _06603_ _02360_ _02362_ _02365_ _02366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12667__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14707_ _01746_ clknet_leaf_88_clk_i memory\[2\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_16_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11919_ _05783_ _06125_ _06127_ _06129_ _06130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_59_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12159__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15687_ _00646_ clknet_leaf_235_clk_i memory\[60\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12899_ _06476_ _02293_ _02295_ _02297_ _02298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__11063__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_99_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14638_ _01677_ clknet_leaf_125_clk_i memory\[27\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_182_clk_i clknet_5_29__leaf_clk_i clknet_leaf_182_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_144_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14569_ _01608_ clknet_leaf_180_clk_i memory\[25\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07110_ _03273_ _00863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08090_ _03831_ _01285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07041_ _03235_ _00832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_197_clk_i clknet_5_28__leaf_clk_i clknet_leaf_197_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_152_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_193_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09261__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12640__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10946__I1 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_120_clk_i clknet_5_23__leaf_clk_i clknet_leaf_120_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08992_ _04325_ _01693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07943_ _03736_ _01233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11238__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07874_ _03194_ memory\[7\]\[22\] _03697_ _03700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09931__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09613_ _04625_ memory\[36\]\[24\] _04664_ _04669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_135_clk_i clknet_5_22__leaf_clk_i clknet_leaf_135_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_108_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_108_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13453__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09544_ _04629_ memory\[35\]\[26\] _04617_ _04630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12577__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07451__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09475_ _03137_ _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__12069__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08426_ _03768_ memory\[20\]\[8\] _04001_ _04010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07250__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08357_ _03973_ _01410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07308_ _03396_ _00938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08282__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08288_ _03766_ memory\[18\]\[7\] _03929_ _03937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07239_ memory\[39\]\[21\] _03353_ _03351_ _03354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11500__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10250_ _05008_ memory\[46\]\[1\] _05006_ _05009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10181_ _04971_ _00156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12532__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09905__I _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07626__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11656__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11148__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_31_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13940_ _00979_ clknet_leaf_130_clk_i memory\[8\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10052__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12934__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_20__f_clk_i clknet_2_2_0_clk_i clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_395_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10987__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13871_ _00910_ clknet_leaf_259_clk_i memory\[39\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15610_ _00569_ clknet_leaf_380_clk_i memory\[57\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12822_ memory\[28\]\[18\] memory\[29\]\[18\] _06604_ _02222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15541_ _00500_ clknet_leaf_42_clk_i memory\[55\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12753_ _02153_ _02154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_29_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11704_ _05681_ _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_16_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10873__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13016__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15472_ _00431_ clknet_leaf_158_clk_i memory\[53\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12684_ _05664_ _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14423_ _01462_ clknet_leaf_98_clk_i memory\[20\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11635_ _05849_ _05850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12707__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11611__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09288__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14354_ _01393_ clknet_leaf_101_clk_i memory\[18\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08192__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09491__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11566_ _05768_ _05771_ _05776_ _05781_ _05782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_141_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13305_ _02367_ _02693_ _02695_ _02697_ _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_162_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10517_ _05041_ memory\[4\]\[17\] _05156_ _05164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14285_ _01324_ clknet_leaf_189_clk_i memory\[29\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11410__I _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11497_ _05710_ _05712_ _05713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13236_ memory\[20\]\[24\] memory\[21\]\[24\] _02368_ _02630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_90_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10448_ _05127_ _00267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13538__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13167_ _02561_ _02562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_104_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10379_ _05039_ memory\[47\]\[16\] _05084_ _05091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11750__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07536__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12118_ _05693_ _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_13098_ _05653_ _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_137_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_52_clk_i clknet_5_18__leaf_clk_i clknet_leaf_52_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12241__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12049_ _05918_ _06257_ _06195_ _06258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07557__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11353__I1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07590_ _03178_ memory\[0\]\[17\] _03541_ _03549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15808_ _00767_ clknet_leaf_301_clk_i memory\[9\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08367__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_67_clk_i clknet_5_16__leaf_clk_i clknet_leaf_67_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15739_ _00698_ clknet_leaf_389_clk_i memory\[61\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13007__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09260_ _04467_ _01819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_103_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08211_ _03896_ _01341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09191_ _04181_ memory\[31\]\[0\] _04430_ _04431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08142_ _03756_ memory\[29\]\[2\] _03857_ _03860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09482__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11664__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08073_ _03822_ _01277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10137__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07024_ net5 _03223_ _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_183_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_140_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10919__I1 _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_149_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11741__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08975_ _04239_ memory\[27\]\[27\] _04308_ _04316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07926_ _03727_ _01225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13494__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input25_I data_i[26] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_162_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07857_ _03169_ memory\[7\]\[14\] _03686_ _03691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_16__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10600__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07788_ _03654_ _01160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_123_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09527_ _04618_ _01935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_151_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09458_ _04571_ _01913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08409_ _04000_ _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09389_ _04245_ memory\[33\]\[30\] _04501_ _04535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12527__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13710__I _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11431__S _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_49_Left_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11420_ _05643_ _00723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09473__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12852__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__I0 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11351_ memory\[61\]\[24\] _03199_ _05602_ _05607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_169_3629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11980__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10302_ _05043_ memory\[46\]\[18\] _05027_ _05044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14070_ _01109_ clknet_leaf_135_clk_i memory\[10\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11282_ _03359_ memory\[60\]\[24\] _05565_ _05570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_186_3943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11032__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13021_ memory\[32\]\[21\] memory\[33\]\[21\] memory\[34\]\[21\] memory\[35\]\[21\]
+ _02205_ _02345_ _02418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12262__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09776__I1 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10233_ _04998_ _00181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07787__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07356__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10164_ _04629_ memory\[44\]\[26\] _04955_ _04962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_58_Left_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14972_ _02011_ clknet_leaf_419_clk_i memory\[38\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10095_ _04925_ _00116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09571__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13923_ _00962_ clknet_leaf_302_clk_i memory\[8\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_141_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11606__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13854_ _00893_ clknet_leaf_418_clk_i memory\[39\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12805_ _05669_ _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13785_ _00824_ clknet_leaf_137_clk_i memory\[14\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10997_ _05043_ memory\[56\]\[18\] _05410_ _05419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15524_ _00483_ clknet_leaf_312_clk_i memory\[55\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10846__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_84_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12736_ _06446_ _02132_ _02134_ _02136_ _02137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_29_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08915__S _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_67_Left_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12945__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_44_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15455_ _00414_ clknet_leaf_331_clk_i memory\[53\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12437__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12667_ _06450_ _06865_ _06866_ _06867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_155_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14406_ _01445_ clknet_leaf_188_clk_i memory\[20\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11618_ _05699_ _05825_ _05832_ _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_61_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09464__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15386_ _00345_ clknet_leaf_380_clk_i memory\[50\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12598_ _06798_ _06799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_142_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14337_ _01376_ clknet_leaf_343_clk_i memory\[18\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11271__I0 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11549_ _05748_ _05751_ _05758_ _05764_ _05765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_41_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11971__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13399__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09216__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14268_ _01307_ clknet_leaf_378_clk_i memory\[29\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_66_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13219_ _02344_ _02612_ _02613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12172__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14199_ _01238_ clknet_leaf_111_clk_i memory\[19\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07778__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07266__S _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Left_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_100_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08760_ _03134_ _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13476__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11326__I1 _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07711_ _03613_ _01124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08691_ _03760_ memory\[24\]\[4\] _04146_ _04151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_68_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10420__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07642_ _03153_ memory\[10\]\[9\] _03567_ _03577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08097__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13228__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07950__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07573_ _03153_ memory\[0\]\[9\] _03530_ _03540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09312_ _04494_ _01844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10837__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07702__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09243_ _04235_ memory\[31\]\[25\] _04452_ _04458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_343_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09174_ _04421_ _01779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09455__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12834__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13400__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08125_ _03849_ _01302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_161_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11962__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09656__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08056_ _03811_ _01271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08560__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09207__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11985__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11014__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07007_ net27 _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_12_672 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput49 net49 data_o[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_164_3526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_164_3537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08958_ _04222_ memory\[27\]\[19\] _04297_ _04307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_181_3851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11317__I1 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09391__S _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07904__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07909_ _03718_ _01217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08889_ _04270_ _01645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08194__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10920_ _05378_ _00488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10330__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09190__I _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10851_ _05341_ _00456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13314__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13570_ _02957_ _02958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08735__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10782_ _05033_ memory\[53\]\[13\] _05301_ _05305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12521_ _06720_ _06722_ _06723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_54_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13078__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15240_ _00199_ clknet_leaf_271_clk_i memory\[46\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12452_ memory\[36\]\[13\] memory\[37\]\[13\] _06447_ _06655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11403_ _05634_ _00715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11253__I0 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15171_ _00130_ clknet_leaf_429_clk_i memory\[44\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12383_ memory\[36\]\[12\] memory\[37\]\[12\] _06447_ _06587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14122_ _01161_ clknet_leaf_224_clk_i memory\[6\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11334_ memory\[61\]\[16\] _03174_ _05591_ _05598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08470__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14053_ _01092_ clknet_leaf_298_clk_i memory\[10\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10505__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11265_ _03342_ memory\[60\]\[16\] _05554_ _05561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07086__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13004_ memory\[6\]\[21\] memory\[7\]\[21\] _02322_ _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10216_ _04989_ _00173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11196_ _05524_ _00618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10304__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10147_ _04612_ memory\[44\]\[18\] _04944_ _04953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07814__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11844__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14955_ _01994_ clknet_leaf_48_clk_i memory\[37\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10078_ _04916_ _00108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_85_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_292_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11564__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11336__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13906_ _00945_ clknet_leaf_120_clk_i memory\[11\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10240__S _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14886_ _01925_ clknet_leaf_48_clk_i memory\[35\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13837_ _00876_ clknet_leaf_195_clk_i memory\[13\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13551__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10819__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13768_ _00807_ clknet_leaf_200_clk_i memory\[14\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09685__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13630__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12719_ memory\[0\]\[17\] memory\[1\]\[17\] memory\[2\]\[17\] memory\[3\]\[17\] _06709_
+ _06779_ _02120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15507_ _00466_ clknet_leaf_154_clk_i memory\[54\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13699_ _03080_ _00767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15438_ _00397_ clknet_leaf_274_clk_i memory\[52\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09437__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12197__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11244__I0 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15369_ _00328_ clknet_leaf_292_clk_i memory\[50\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11944__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12292__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09476__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09930_ _04838_ _00038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Right_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_159_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09861_ _04598_ memory\[40\]\[11\] _04800_ _04802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08812_ _03186_ _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_142_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09792_ _04764_ _02054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13449__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08743_ _03812_ memory\[24\]\[29\] _04168_ _04178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11246__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12121__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08674_ _04141_ _01559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07923__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_96_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_120_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07625_ _03568_ _01083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_24_Right_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_193_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_113_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07556_ _03531_ _01051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13621__A1 _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12585__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07487_ _03494_ _01019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09226_ _04218_ memory\[31\]\[17\] _04441_ _04449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09428__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_118_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_118_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09157_ _04412_ _01771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08108_ _03840_ _01294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_135_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08290__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09088_ _04216_ memory\[2\]\[16\] _04369_ _04376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_169_Right_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_163_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_33_Right_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_130_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08039_ _03196_ _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_3_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_183_3902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12035__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11050_ _05447_ _00549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09600__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10001_ _04602_ memory\[42\]\[13\] _04872_ _04876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12540__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output56_I net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08167__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14740_ _01779_ clknet_leaf_90_clk_i memory\[30\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10060__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11952_ _05667_ _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_19_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07914__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_42_Right_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10903_ _05369_ _00480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14671_ _01710_ clknet_leaf_183_clk_i memory\[28\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10995__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_28_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11883_ memory\[12\]\[5\] memory\[13\]\[5\] _06025_ _06094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13371__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13622_ _02964_ _02979_ _02994_ _03009_ _03010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_10834_ _05332_ _00448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13612__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13553_ memory\[22\]\[29\] memory\[23\]\[29\] _05754_ _02942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10765_ _05016_ memory\[53\]\[5\] _05290_ _05296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12504_ memory\[6\]\[14\] memory\[7\]\[14\] _06431_ _06706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13484_ _02498_ _02873_ _05665_ _02874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10696_ _05259_ _00383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11226__I0 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15223_ _00182_ clknet_leaf_17_clk_i memory\[45\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_239_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12435_ _06142_ _06633_ _06635_ _06637_ _06638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_113_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12715__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_51_Right_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09296__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15154_ _00113_ clknet_leaf_13_clk_i memory\[43\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12366_ _06411_ _06562_ _06569_ _06570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08642__I1 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_136_Right_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14105_ _01144_ clknet_leaf_146_clk_i memory\[63\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11317_ memory\[61\]\[8\] _03149_ _05580_ _05589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_39_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15085_ _00044_ clknet_leaf_23_clk_i memory\[41\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12297_ memory\[54\]\[11\] memory\[55\]\[11\] _06421_ _06502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14036_ _01075_ clknet_leaf_57_clk_i memory\[0\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11248_ _03325_ memory\[60\]\[8\] _05543_ _05552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_56_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13546__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11179_ _05515_ _00610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07544__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_60_Right_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14938_ _01977_ clknet_leaf_444_clk_i memory\[36\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07343__I _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14869_ _01908_ clknet_leaf_74_clk_i memory\[34\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07410_ net5 net6 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08375__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08390_ _03800_ memory\[1\]\[23\] _03987_ _03991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09658__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07341_ _03413_ _00954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08330__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07272_ _03265_ _03375_ _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
Xclkbuf_leaf_411_clk_i clknet_5_2__leaf_clk_i clknet_leaf_411_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_14_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09011_ _04335_ _01702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_72_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12625__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13462__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07719__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08633__I1 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_76_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_103_Right_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_426_clk_i clknet_5_0__leaf_clk_i clknet_leaf_426_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10145__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09913_ _04829_ _00030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_130_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09844_ _04581_ memory\[40\]\[3\] _04789_ _04793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09775_ _04755_ _02046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06987_ net22 _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11528__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08726_ _04169_ _01583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08849__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07253__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_188_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08657_ memory\[23\]\[20\] _03350_ _04132_ _04133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_159_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13191__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07608_ _03558_ _01076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08588_ _03793_ memory\[22\]\[20\] _04095_ _04096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09649__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_176_3761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_36_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07539_ _03521_ _01044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11503__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10550_ _05004_ memory\[50\]\[0\] _05181_ _05182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_240_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11208__I0 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09209_ _04201_ memory\[31\]\[9\] _04430_ _04440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10481_ _05144_ _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_161_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12220_ _06142_ _06420_ _06423_ _06425_ _06426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08812__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11659__B _05870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12581__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12151_ memory\[54\]\[9\] memory\[55\]\[9\] _05684_ _06358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11102_ _03315_ memory\[58\]\[3\] _05471_ _05475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09844__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12082_ _06149_ _06289_ _06290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08388__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_21_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11033_ _05438_ _00541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15772_ _00731_ clknet_leaf_349_clk_i net40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09888__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12984_ _03122_ _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_87_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14723_ _01762_ clknet_leaf_409_clk_i memory\[30\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11935_ _06144_ _06145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08560__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14654_ _01693_ clknet_leaf_354_clk_i memory\[28\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11866_ _05654_ _06072_ _06074_ _06076_ _06077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_28_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13605_ _05676_ _02988_ _02990_ _02992_ _02993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10817_ _05068_ memory\[53\]\[30\] _05289_ _05323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14585_ _01624_ clknet_leaf_78_clk_i memory\[25\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11797_ _05682_ _06008_ _05687_ _06009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_131_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13536_ memory\[44\]\[29\] memory\[45\]\[29\] _05678_ _02925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08923__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10748_ _05286_ _00408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_164_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13467_ _02856_ _02857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_97_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10679_ memory\[51\]\[29\] _03214_ _05240_ _05250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15206_ _00165_ clknet_leaf_32_clk_i memory\[45\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12418_ _06467_ _06614_ _06621_ _06622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_23_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13398_ _05772_ _02788_ _02195_ _02789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08615__I1 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12572__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15137_ _00096_ clknet_leaf_439_clk_i memory\[43\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12349_ _06553_ net42 _06491_ _06554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12244__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15068_ _00027_ clknet_leaf_434_clk_i memory\[41\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08379__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_442_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14019_ _01058_ clknet_leaf_336_clk_i memory\[0\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06910_ _03137_ _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_103_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10186__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07890_ _03218_ memory\[7\]\[30\] _03674_ _03708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_71_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07051__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11922__I1 net67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09560_ _04640_ _01946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08511_ _03785_ memory\[21\]\[16\] _04048_ _04055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12183__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09491_ _04593_ memory\[35\]\[9\] _04575_ _04594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_19_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08442_ _04018_ _01450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_19_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07801__I _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_137_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08373_ _03783_ memory\[1\]\[15\] _03976_ _03982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08303__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_350_clk_i clknet_5_8__leaf_clk_i clknet_leaf_350_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07324_ memory\[11\]\[23\] _03357_ _03401_ _03405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_154_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09929__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10110__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_12_Left_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_116_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_469 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07255_ _03364_ _00917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_115_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10661__I1 _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07449__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_365_clk_i clknet_5_9__leaf_clk_i clknet_leaf_365_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07186_ memory\[39\]\[4\] _03317_ _03309_ _03318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09664__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12315__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13186__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11749__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_21_Left_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09463__I _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07042__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09827_ _04782_ _02071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09758_ _04745_ _02039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_303_clk_i clknet_5_14__leaf_clk_i clknet_leaf_303_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_178_3801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07912__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08709_ _04160_ _01575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09689_ _04633_ memory\[37\]\[28\] _04700_ _04709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08542__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11720_ _05881_ _05897_ _05913_ _05933_ _05934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_51_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11429__I0 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11651_ _05865_ _00732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_318_clk_i clknet_5_11__leaf_clk_i clknet_leaf_318_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_30_Left_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_181_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13674__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_10602_ _05058_ memory\[50\]\[25\] _05203_ _05209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14370_ _01409_ clknet_leaf_339_clk_i memory\[1\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08743__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11582_ _05794_ _05797_ _05798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_391_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13321_ memory\[48\]\[26\] memory\[49\]\[26\] memory\[50\]\[26\] memory\[51\]\[26\]
+ _05725_ _05726_ _02713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_107_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10533_ _05172_ _00307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__I1 _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13252_ _02170_ _02644_ _02645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10464_ _05056_ memory\[48\]\[24\] _05131_ _05136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12203_ _06409_ net71 _05802_ _06410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12064__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13183_ _02577_ _00754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_5__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10395_ _05099_ _00242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12134_ _05691_ _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_20_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12306__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12065_ _05655_ _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10513__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10168__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07094__S _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11016_ _05062_ memory\[56\]\[27\] _05421_ _05429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15824_ _00783_ clknet_leaf_126_clk_i memory\[9\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07822__S _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11852__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12967_ _06610_ _02364_ _02365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15755_ _00714_ clknet_leaf_225_clk_i memory\[62\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07336__I1 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14706_ _01745_ clknet_leaf_58_clk_i memory\[2\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11918_ _05794_ _06128_ _06129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_34_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_16_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12898_ _06484_ _02296_ _02297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15686_ _00645_ clknet_leaf_236_clk_i memory\[60\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14637_ _01676_ clknet_leaf_124_clk_i memory\[27\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11849_ _06060_ _06061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12239__I _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09749__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14568_ _01607_ clknet_leaf_183_clk_i memory\[25\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13519_ _05759_ _02907_ _02908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14499_ _01538_ clknet_leaf_356_clk_i memory\[23\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07269__S _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07040_ _03141_ memory\[16\]\[5\] _03229_ _03235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_136_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12545__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12640__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08991_ _04187_ memory\[28\]\[2\] _04322_ _04325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_76_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07942_ _03194_ memory\[19\]\[22\] _03733_ _03736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07873_ _03699_ _01200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13734__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09612_ _04668_ _01970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_108_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_108_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09543_ _03205_ _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08524__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12320__I1 memory\[39\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09474_ _04582_ _01918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_38_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08425_ _04009_ _01442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08356_ _03766_ memory\[1\]\[7\] _03965_ _03973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12593__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07307_ memory\[11\]\[15\] _03340_ _03390_ _03396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08287_ _03936_ _01377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12085__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08362__I _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07238_ _03190_ _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_132_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08204__A2 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07169_ _03112_ _03304_ _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10398__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10180_ _04577_ memory\[45\]\[1\] _04969_ _04971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11429__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10333__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_338_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12395__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_31_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_242_clk_i clknet_5_26__leaf_clk_i clknet_leaf_242_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13870_ _00909_ clknet_leaf_259_clk_i memory\[39\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07642__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12821_ _06445_ _02208_ _02220_ _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08515__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07318__I1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12752_ memory\[20\]\[17\] memory\[21\]\[17\] _06477_ _02153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15540_ _00499_ clknet_leaf_154_clk_i memory\[55\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_257_clk_i clknet_5_13__leaf_clk_i clknet_leaf_257_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_16_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11703_ _05916_ _05917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_166_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15471_ _00430_ clknet_leaf_274_clk_i memory\[53\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12683_ memory\[30\]\[16\] memory\[31\]\[16\] _02084_ _02085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14422_ _01461_ clknet_leaf_93_clk_i memory\[20\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09569__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11634_ memory\[28\]\[1\] memory\[29\]\[1\] _05769_ _05849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_46_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14353_ _01392_ clknet_leaf_102_clk_i memory\[18\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10625__I1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11565_ _05777_ _05780_ _05781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_107_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13304_ _02375_ _02696_ _02697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09368__I _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10516_ _05163_ _00299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14284_ _01323_ clknet_leaf_184_clk_i memory\[29\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11496_ memory\[0\]\[0\] memory\[1\]\[0\] memory\[2\]\[0\] memory\[3\]\[0\] _05711_
+ _03748_ _05712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_134_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13235_ _02494_ _02624_ _02626_ _02628_ _02629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10307__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10447_ _05039_ memory\[48\]\[16\] _05120_ _05127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13166_ memory\[28\]\[23\] memory\[29\]\[23\] _02495_ _02561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10378_ _05090_ _00234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11750__A2 _05962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12117_ _05689_ _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_13097_ _02336_ _02484_ _02492_ _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_100_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12048_ memory\[30\]\[7\] memory\[31\]\[7\] _06193_ _06257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15807_ _00766_ clknet_leaf_309_clk_i memory\[9\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07309__I1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11074__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13999_ _01038_ clknet_leaf_242_clk_i memory\[59\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_62_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15738_ _00697_ clknet_leaf_388_clk_i memory\[61\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_190_4020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15669_ _00628_ clknet_leaf_142_clk_i memory\[5\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08210_ _03756_ memory\[17\]\[2\] _03893_ _03896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_83_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09479__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09190_ _04429_ _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13558__A3 _02946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08141_ _03859_ _01308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13302__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10418__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08072_ _03756_ memory\[15\]\[2\] _03819_ _03822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_287_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13729__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07023_ net6 _03223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_2
XFILLER_0_12_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12633__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07727__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08993__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11741__A2 _05953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08974_ _04315_ _01685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_89_Right_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07925_ _03169_ memory\[19\]\[14\] _03722_ _03727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11048__I _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08745__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07548__I1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07856_ _03690_ _01192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_162_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08558__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10552__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07462__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input18_I data_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07787_ _03166_ memory\[6\]\[13\] _03650_ _03654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_123_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_123_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09526_ _04616_ memory\[35\]\[20\] _04617_ _04618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_79_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09457_ _04245_ memory\[34\]\[30\] _04537_ _04571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13629__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11712__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09389__S _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08408_ _03225_ _03750_ _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XPHY_EDGE_ROW_98_Right_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10480__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09388_ _04534_ _01880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08339_ _03963_ _01402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12852__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12221__A3 _06426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11350_ _05606_ _00690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12509__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10301_ _03180_ _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_132_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11281_ _05569_ _00658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13020_ _02341_ _02416_ _06866_ _02417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_186_3944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10232_ _04629_ memory\[45\]\[26\] _04991_ _04998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_186_3955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10063__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10163_ _04961_ _00148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_5_Left_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_7_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_181_clk_i clknet_5_28__leaf_clk_i clknet_leaf_181_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09852__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07436__I _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14971_ _02010_ clknet_leaf_443_clk_i memory\[37\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10094_ _04627_ memory\[43\]\[25\] _04919_ _04925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13922_ _00961_ clknet_leaf_302_clk_i memory\[8\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08468__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09651__I _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13853_ _00892_ clknet_leaf_411_clk_i memory\[39\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_196_clk_i clknet_5_29__leaf_clk_i clknet_leaf_196_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_186_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_48_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12804_ _06450_ _02203_ _06866_ _02204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13784_ _00823_ clknet_leaf_140_clk_i memory\[14\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10996_ _05418_ _00524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15523_ _00482_ clknet_leaf_335_clk_i memory\[55\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12735_ _06453_ _02135_ _02136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_44_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15454_ _00413_ clknet_leaf_346_clk_i memory\[53\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12666_ _05686_ _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12748__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14405_ _01444_ clknet_leaf_375_clk_i memory\[20\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11617_ _05715_ _05827_ _05829_ _05831_ _05832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_53_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_61_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10238__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15385_ _00344_ clknet_leaf_381_clk_i memory\[50\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12597_ memory\[44\]\[15\] memory\[45\]\[15\] _06319_ _06798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14336_ _01375_ clknet_leaf_348_clk_i memory\[18\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11548_ _05760_ _05763_ _05764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08931__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_134_clk_i clknet_5_22__leaf_clk_i clknet_leaf_134_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_40_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14267_ _01306_ clknet_leaf_394_clk_i memory\[15\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11479_ memory\[48\]\[0\] memory\[49\]\[0\] memory\[50\]\[0\] memory\[51\]\[0\] _05692_
+ _05694_ _05695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_64_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13218_ memory\[32\]\[24\] memory\[33\]\[24\] memory\[34\]\[24\] memory\[35\]\[24\]
+ _02205_ _02345_ _02612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11577__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14198_ _01237_ clknet_leaf_110_clk_i memory\[19\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12920__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08975__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13149_ _06713_ _02539_ _02541_ _02543_ _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_0_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_149_clk_i clknet_5_19__leaf_clk_i clknet_leaf_149_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10782__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08727__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13284__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07710_ _03153_ memory\[63\]\[9\] _03603_ _03613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_144_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10701__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08690_ _04150_ _01566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10534__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07282__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07641_ _03576_ _01091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_105_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07572_ _03539_ _01059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09152__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09311_ _04235_ memory\[32\]\[25\] _04488_ _04494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_165_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09242_ _04457_ _01811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09173_ _04233_ memory\[30\]\[24\] _04416_ _04421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_111_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12834__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08124_ _03808_ memory\[15\]\[27\] _03841_ _03849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09937__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08841__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08055_ _03810_ memory\[12\]\[28\] _03794_ _03811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07006_ _03210_ _00822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13164__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12911__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_164_3538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10773__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07256__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08957_ _04306_ _01677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_181_3863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08718__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13711__I0 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07908_ _03144_ memory\[19\]\[6\] _03711_ _03718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08888_ _04220_ memory\[26\]\[18\] _04261_ _04270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08288__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07192__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09391__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07839_ _03681_ _01184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11506__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10850_ _05033_ memory\[54\]\[13\] _05337_ _05341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09509_ _03171_ _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10781_ _05304_ _00423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12520_ memory\[8\]\[14\] memory\[9\]\[14\] memory\[10\]\[14\] memory\[11\]\[14\]
+ _06582_ _06721_ _06722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_137_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_93_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13078__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_117_Right_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_23_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12451_ _06428_ _06646_ _06653_ _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__10058__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_51_clk_i clknet_5_19__leaf_clk_i clknet_leaf_51_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_164_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11402_ _03342_ memory\[62\]\[16\] _05627_ _05634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15170_ _00129_ clknet_leaf_432_clk_i memory\[44\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12382_ _06428_ _06577_ _06585_ _06586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_14121_ _01160_ clknet_leaf_223_clk_i memory\[6\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_10_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11333_ _05597_ _00682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07367__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14052_ _01091_ clknet_leaf_294_clk_i memory\[10\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_66_clk_i clknet_5_16__leaf_clk_i clknet_leaf_66_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11264_ _05560_ _00650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13003_ _02399_ _02400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_120_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12072__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10215_ _04612_ memory\[45\]\[18\] _04980_ _04989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11195_ _03340_ memory\[5\]\[15\] _05518_ _05524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10146_ _04952_ _00140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13702__I0 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10521__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08198__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10077_ _04610_ memory\[43\]\[17\] _04908_ _04916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14954_ _01993_ clknet_leaf_49_clk_i memory\[37\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_235_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13905_ _00944_ clknet_leaf_121_clk_i memory\[11\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11564__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_85_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14885_ _01924_ clknet_leaf_400_clk_i memory\[35\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10320__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13836_ _00875_ clknet_leaf_198_clk_i memory\[13\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07830__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_174_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13767_ _00806_ clknet_leaf_218_clk_i memory\[14\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10979_ _05409_ _00516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09834__A1 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15506_ _00465_ clknet_leaf_154_clk_i memory\[54\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12718_ _06848_ _02118_ _06707_ _02119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07696__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13698_ _03317_ memory\[9\]\[4\] _03075_ _03080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_19_clk_i clknet_5_5__leaf_clk_i clknet_leaf_19_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15437_ _00396_ clknet_leaf_289_clk_i memory\[52\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12247__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12649_ memory\[6\]\[16\] memory\[7\]\[16\] _06431_ _06849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13394__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09757__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08661__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15368_ _00327_ clknet_leaf_292_clk_i memory\[50\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13279__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14319_ _01358_ clknet_leaf_193_clk_i memory\[17\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15299_ _00258_ clknet_leaf_315_clk_i memory\[48\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13146__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08948__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09860_ _04801_ _00005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10755__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08811_ _04223_ _01614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09791_ memory\[3\]\[11\] _03159_ _04762_ _04764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08742_ _04177_ _01591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10507__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09373__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08673_ memory\[23\]\[28\] _03367_ _04132_ _04141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13027__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11180__I0 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13742__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07624_ _03111_ memory\[10\]\[0\] _03567_ _03568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_120_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12866__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07740__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09125__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07555_ _03111_ memory\[0\]\[0\] _03530_ _03531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_75_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11632__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_437_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08635__I _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07486_ memory\[59\]\[0\] _03303_ _03493_ _03494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09225_ _04448_ _01803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_157_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_8_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13385__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09156_ _04216_ memory\[30\]\[16\] _04405_ _04412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08571__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_118_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09053__A2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08107_ _03791_ memory\[15\]\[19\] _03830_ _03840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09087_ _04375_ _01738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_135_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10606__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_184_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09466__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08038_ _03799_ _01265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_3903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13688__A2 net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11699__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10000_ _04875_ _00071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07611__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12991__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09989_ _04869_ _00066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09364__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output49_I net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_95_Left_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11951_ _06159_ _06160_ _06018_ _06161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_99_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_28_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10902_ memory\[55\]\[5\] _03140_ _05363_ _05369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14670_ _01709_ clknet_leaf_183_clk_i memory\[28\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_28_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11882_ _05700_ _06087_ _06089_ _06092_ _06093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_54_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10833_ _05016_ memory\[54\]\[5\] _05326_ _05332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13621_ _03224_ _03001_ _03008_ _03009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_67_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11172__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07678__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13552_ _02940_ _02941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10764_ _05295_ _00415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08545__I _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12503_ _06704_ _06705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13483_ memory\[30\]\[28\] memory\[31\]\[28\] _05737_ _02873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10695_ _05014_ memory\[52\]\[4\] _05254_ _05259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13376__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11900__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09577__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15222_ _00181_ clknet_leaf_15_clk_i memory\[45\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12434_ _06149_ _06636_ _06637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15153_ _00112_ clknet_leaf_8_clk_i memory\[43\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12365_ _06142_ _06564_ _06566_ _06568_ _06569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__10985__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14104_ _01143_ clknet_leaf_145_clk_i memory\[63\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11316_ _05588_ _00674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_22_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15084_ _00043_ clknet_leaf_25_clk_i memory\[41\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12296_ _06500_ _06501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_39_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14035_ _01074_ clknet_leaf_139_clk_i memory\[0\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11247_ _05551_ _00642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_56_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10737__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11178_ _03323_ memory\[5\]\[7\] _05507_ _05515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11347__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10129_ _04943_ _00132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_386_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12734__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14937_ _01976_ clknet_leaf_14_clk_i memory\[36\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13562__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14868_ _01907_ clknet_leaf_74_clk_i memory\[34\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13819_ _00858_ clknet_leaf_28_clk_i memory\[16\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14799_ _01838_ clknet_leaf_51_clk_i memory\[32\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11082__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07340_ memory\[11\]\[31\] _03373_ _03378_ _03413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_139_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11614__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07271_ _03116_ _03264_ _03375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_0_45_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09010_ _04206_ memory\[28\]\[11\] _04333_ _04335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13367__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13462__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10426__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10976__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09830__I1 _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09912_ _04581_ memory\[41\]\[3\] _04825_ _04829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09594__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09843_ _04792_ _02077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11257__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06986_ _03195_ _00817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09774_ memory\[3\]\[3\] _03134_ _04751_ _04755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09950__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11528__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08725_ _03793_ memory\[24\]\[20\] _04168_ _04169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08656_ _04109_ _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07470__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07607_ _03203_ memory\[0\]\[25\] _03552_ _03558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_159_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08587_ _04072_ _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_49_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07538_ memory\[59\]\[25\] _03361_ _03515_ _03521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_14_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07469_ _03483_ _01012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13358__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09208_ _04439_ _01795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10480_ _03528_ _03750_ _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_17_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09139_ _04199_ memory\[30\]\[8\] _04394_ _04403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12030__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10336__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_14__f_clk_i clknet_2_1_0_clk_i clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_121_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12581__A2 _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12150_ _06356_ _06357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07832__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11101_ _05474_ _00573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13647__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12081_ memory\[48\]\[8\] memory\[49\]\[8\] memory\[50\]\[8\] memory\[51\]\[8\] _06010_
+ _06150_ _06289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_25_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07645__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11032_ _05010_ memory\[57\]\[2\] _05435_ _05438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10344__A1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11392__I0 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_34_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_34_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10071__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09337__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12097__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15771_ _00730_ clknet_leaf_389_clk_i memory\[62\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12983_ _02318_ _02335_ _02357_ _02380_ _02381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__11144__I0 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13382__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14722_ _01761_ clknet_leaf_410_clk_i memory\[30\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11844__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11934_ memory\[52\]\[6\] memory\[53\]\[6\] _06143_ _06144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_170_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14653_ _01692_ clknet_leaf_389_clk_i memory\[28\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11865_ _05668_ _06075_ _06076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_32_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13604_ _05690_ _02991_ _02992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__13597__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10816_ _05322_ _00440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14584_ _01623_ clknet_leaf_78_clk_i memory\[25\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11796_ memory\[54\]\[4\] memory\[55\]\[4\] _05684_ _06008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13535_ _02337_ _02919_ _02921_ _02923_ _02924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_54_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10747_ _05066_ memory\[52\]\[29\] _05276_ _05286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10678_ _05249_ _00375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13466_ memory\[36\]\[28\] memory\[37\]\[28\] _02338_ _02856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_97_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15205_ _00164_ clknet_leaf_430_clk_i memory\[45\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12417_ _06476_ _06616_ _06618_ _06620_ _06621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_153_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12021__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08076__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13397_ memory\[14\]\[27\] memory\[15\]\[27\] _02193_ _02788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_58_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09812__I1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15136_ _00095_ clknet_leaf_439_clk_i memory\[43\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12348_ _06507_ _06522_ _06537_ _06552_ _06553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_12279_ _05693_ _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_15067_ _00026_ clknet_leaf_443_clk_i memory\[40\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12461__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07555__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12324__A2 _06524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14018_ _01057_ clknet_leaf_337_clk_i memory\[0\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11383__I0 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09770__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12088__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11135__I0 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_132_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08510_ _04054_ _01482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13292__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11805__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08000__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12183__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09490_ _03152_ _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_188_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08386__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08441_ _03783_ memory\[20\]\[15\] _04012_ _04018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13091__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13132__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08372_ _03981_ _01417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_193_4095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07323_ _03404_ _00945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12260__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12636__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07254_ memory\[39\]\[26\] _03363_ _03351_ _03364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_115_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09010__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_30_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07185_ _03137_ _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10156__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09803__I1 _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_132_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07814__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09945__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_57_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07290__I1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09567__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13512__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11749__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09826_ memory\[3\]\[28\] _03211_ _04773_ _04782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09319__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09757_ _04633_ memory\[38\]\[28\] _04736_ _04745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06969_ _03182_ _00813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08708_ _03777_ memory\[24\]\[12\] _04157_ _04160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09688_ _04708_ _02006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_169_Left_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_68_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08639_ _04123_ _01542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11650_ _05864_ net51 _05802_ _05865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13674__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10601_ _05208_ _00339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11581_ memory\[16\]\[0\] memory\[17\]\[0\] memory\[18\]\[0\] memory\[19\]\[0\] _05795_
+ _05796_ _05797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_65_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_334_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10532_ _05056_ memory\[4\]\[24\] _05167_ _05172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13320_ _05719_ _02711_ _02178_ _02712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_51_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08058__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13251_ memory\[56\]\[25\] memory\[57\]\[25\] memory\[58\]\[25\] memory\[59\]\[25\]
+ _06827_ _02171_ _02644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10463_ _05135_ _00274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_162_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_178_Left_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12202_ _06363_ _06378_ _06393_ _06408_ _06409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_13182_ _02576_ net55 _02382_ _02577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10394_ _05054_ memory\[47\]\[23\] _05095_ _05099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_92_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12133_ _05788_ _06340_ _05792_ _06341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_92_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07375__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12064_ _05653_ _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_11015_ _05428_ _00533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_410_clk_i clknet_5_2__leaf_clk_i clknet_leaf_410_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09590__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15823_ _00782_ clknet_leaf_203_clk_i memory\[9\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11117__I0 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_187_Left_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15754_ _00713_ clknet_leaf_225_clk_i memory\[62\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12966_ memory\[24\]\[20\] memory\[25\]\[20\] memory\[26\]\[20\] memory\[27\]\[20\]
+ _02363_ _06611_ _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_73_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14705_ _01744_ clknet_leaf_89_clk_i memory\[2\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09730__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11917_ memory\[16\]\[5\] memory\[17\]\[5\] memory\[18\]\[5\] memory\[19\]\[5\] _05795_
+ _05796_ _06128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_87_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15685_ _00644_ clknet_leaf_306_clk_i memory\[60\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12897_ memory\[16\]\[19\] memory\[17\]\[19\] memory\[18\]\[19\] memory\[19\]\[19\]
+ _02233_ _06485_ _02296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_16_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_425_clk_i clknet_5_0__leaf_clk_i clknet_leaf_425_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13114__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14636_ _01675_ clknet_leaf_186_clk_i memory\[27\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11848_ memory\[20\]\[4\] memory\[21\]\[4\] _05785_ _06060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12964__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08297__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14567_ _01606_ clknet_leaf_178_clk_i memory\[25\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11779_ memory\[16\]\[3\] memory\[17\]\[3\] memory\[18\]\[3\] memory\[19\]\[3\] _05795_
+ _05796_ _05992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_166_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13518_ memory\[0\]\[29\] memory\[1\]\[29\] memory\[2\]\[29\] memory\[3\]\[29\] _05784_
+ _03226_ _02907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_14498_ _01537_ clknet_leaf_358_clk_i memory\[23\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_82_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_841 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08049__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12255__I _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13449_ _05715_ _02834_ _02836_ _02838_ _02839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_2_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15119_ _00078_ clknet_leaf_19_clk_i memory\[42\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08990_ _04324_ _01692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07941_ _03735_ _01232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07872_ _03191_ memory\[7\]\[21\] _03697_ _03699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11600__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09611_ _04623_ memory\[36\]\[23\] _04664_ _04668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11108__I0 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_283_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_108_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_108_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09542_ _04628_ _01940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_125_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09005__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13035__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12481__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09473_ _04581_ memory\[35\]\[3\] _04575_ _04582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13750__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08424_ _03766_ memory\[20\]\[7\] _04001_ _04009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08844__S _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12874__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08288__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08355_ _03972_ _01409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07306_ _03395_ _00937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08286_ _03764_ memory\[18\]\[6\] _03929_ _03936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07237_ _03352_ _00911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09675__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07259__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07168_ net5 _03223_ _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__or2_4
XANTENNA__07412__A1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08460__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07263__I1 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10614__S _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07099_ _03115_ net76 _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_100_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07195__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11509__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08212__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10413__I _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12395__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07923__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09960__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09809_ _04750_ _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_92_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12820_ _02209_ _02212_ _02215_ _02219_ _02220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__13344__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12751_ _06603_ _02147_ _02149_ _02151_ _02152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12472__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11702_ memory\[28\]\[2\] memory\[29\]\[2\] _05915_ _05916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15470_ _00429_ clknet_leaf_274_clk_i memory\[53\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12682_ _05683_ _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_167_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13016__A3 _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14421_ _01460_ clknet_leaf_100_clk_i memory\[20\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_127_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11633_ _05731_ _05840_ _05847_ _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_181_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11180__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10086__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14352_ _01391_ clknet_leaf_103_clk_i memory\[18\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11564_ memory\[24\]\[0\] memory\[25\]\[0\] memory\[26\]\[0\] memory\[27\]\[0\] _05778_
+ _05779_ _05780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_64_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13303_ memory\[16\]\[25\] memory\[17\]\[25\] memory\[18\]\[25\] memory\[19\]\[25\]
+ _02233_ _02376_ _02696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_94_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10515_ _05039_ memory\[4\]\[16\] _05156_ _05163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14283_ _01322_ clknet_leaf_188_clk_i memory\[29\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11495_ _03120_ _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13234_ _02501_ _02627_ _02628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10446_ _05126_ _00266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_90_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_110_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15585__CLK clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10524__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10377_ _05037_ memory\[47\]\[15\] _05084_ _05090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07254__I1 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13165_ _02336_ _02552_ _02559_ _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__11830__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12116_ _06322_ _06323_ _05757_ _06324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13096_ _02209_ _02486_ _02489_ _02491_ _02492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_104_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12047_ _06255_ _06256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10323__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08929__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11863__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11355__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15806_ _00765_ clknet_leaf_309_clk_i memory\[9\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13998_ _01037_ clknet_leaf_243_clk_i memory\[59\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09703__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_364_clk_i clknet_5_9__leaf_clk_i clknet_leaf_364_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_62_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15737_ _00696_ clknet_leaf_382_clk_i memory\[61\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12949_ _02344_ _02346_ _02347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_158_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_29_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_66_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_66_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_190_4021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15668_ _00627_ clknet_leaf_142_clk_i memory\[5\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_103_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_29_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14619_ _01658_ clknet_leaf_5_clk_i memory\[26\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15599_ _00558_ clknet_leaf_243_clk_i memory\[57\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_379_clk_i clknet_5_12__leaf_clk_i clknet_leaf_379_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11090__S _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08140_ _03754_ memory\[29\]\[1\] _03857_ _03859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10077__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08071_ _03821_ _01276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07022_ _03222_ _00826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09495__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_302_clk_i clknet_5_14__leaf_clk_i clknet_leaf_302_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_141_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__I1 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11821__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_149_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_149_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08973_ _04237_ memory\[27\]\[26\] _04308_ _04315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_317_clk_i clknet_5_11__leaf_clk_i clknet_leaf_317_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_166_3580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07924_ _03726_ _01224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10001__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07855_ _03166_ memory\[7\]\[13\] _03686_ _03690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_162_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11265__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07786_ _03653_ _01159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09525_ _04574_ _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_52_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09456_ _04570_ _01912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13629__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08407_ _03999_ _01434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_191_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09387_ _04243_ memory\[33\]\[29\] _04524_ _04534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09469__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12757__A2 _02157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08338_ _03816_ memory\[18\]\[31\] _03928_ _03963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08269_ _03926_ _01369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12824__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10300_ _05042_ _00204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11280_ _03357_ memory\[60\]\[23\] _05565_ _05569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10231_ _04997_ _00180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_186_3945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08433__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07236__I1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10240__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10162_ _04627_ memory\[44\]\[25\] _04955_ _04961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13655__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14970_ _02009_ clknet_leaf_443_clk_i memory\[37\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10093_ _04924_ _00115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07653__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12779__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09933__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13921_ _00960_ clknet_leaf_301_clk_i memory\[8\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13852_ _00891_ clknet_leaf_411_clk_i memory\[39\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_87_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_179_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12803_ memory\[38\]\[18\] memory\[39\]\[18\] _06728_ _02203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13783_ _00822_ clknet_leaf_135_clk_i memory\[14\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10995_ _05041_ memory\[56\]\[17\] _05410_ _05418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13390__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15522_ _00481_ clknet_leaf_335_clk_i memory\[55\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12734_ memory\[32\]\[17\] memory\[33\]\[17\] memory\[34\]\[17\] memory\[35\]\[17\]
+ _06314_ _06454_ _02135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_123_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08484__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15453_ _00412_ clknet_leaf_345_clk_i memory\[53\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10519__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12665_ memory\[38\]\[16\] memory\[39\]\[16\] _06728_ _06865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14404_ _01443_ clknet_leaf_377_clk_i memory\[20\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11616_ _05724_ _05830_ _05831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_61_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15384_ _00343_ clknet_leaf_381_clk_i memory\[50\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12596_ _06446_ _06792_ _06794_ _06796_ _06797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_61_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12019__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_231_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14335_ _01374_ clknet_leaf_356_clk_i memory\[18\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11547_ memory\[40\]\[0\] memory\[41\]\[0\] memory\[42\]\[0\] memory\[43\]\[0\] _05761_
+ _05762_ _05763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_123_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07828__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14266_ _01305_ clknet_leaf_31_clk_i memory\[15\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11478_ _05693_ _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13217_ _02341_ _02610_ _06866_ _02611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10429_ _05117_ _00258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08424__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14197_ _01236_ clknet_leaf_115_clk_i memory\[19\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13148_ _06720_ _02542_ _02543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13079_ _06720_ _02474_ _02475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08659__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07563__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09924__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_68_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07640_ _03150_ memory\[10\]\[8\] _03567_ _03576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_105_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13228__A3 _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07571_ _03150_ memory\[0\]\[8\] _03530_ _03539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12436__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09310_ _04493_ _01843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08394__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06907__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07163__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09241_ _04233_ memory\[31\]\[24\] _04452_ _04457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13313__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09172_ _04420_ _01778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08123_ _03848_ _01301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_241_clk_i clknet_5_13__leaf_clk_i clknet_leaf_241_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07466__I1 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07738__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08054_ _03211_ _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10470__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07005_ _03209_ memory\[14\]\[27\] _03188_ _03210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10164__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10222__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_256_clk_i clknet_5_24__leaf_clk_i clknet_leaf_256_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06977__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_164_3539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_433_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13475__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08956_ _04220_ memory\[27\]\[18\] _04297_ _04306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08569__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input30_I data_i[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07907_ _03717_ _01216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08887_ _04269_ _01644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07838_ _03141_ memory\[7\]\[5\] _03675_ _03681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_180_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12427__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07769_ _03644_ _01151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11723__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09508_ _04605_ _01929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10780_ _05031_ memory\[53\]\[12\] _05301_ _05304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09439_ _04227_ memory\[34\]\[21\] _04560_ _04562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10339__S _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12450_ _06024_ _06648_ _06650_ _06652_ _06653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_23_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_209_clk_i clknet_5_30__leaf_clk_i clknet_leaf_209_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_191_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11401_ _05633_ _00714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12381_ _06024_ _06579_ _06581_ _06584_ _06585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_105_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14120_ _01159_ clknet_leaf_222_clk_i memory\[6\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08831__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11332_ memory\[61\]\[15\] _03171_ _05591_ _05597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11678__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12353__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08406__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14051_ _01090_ clknet_leaf_301_clk_i memory\[10\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11263_ _03340_ memory\[60\]\[15\] _05554_ _05560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13002_ memory\[4\]\[21\] memory\[5\]\[21\] _06845_ _02399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09863__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10213__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10214_ _04988_ _00172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11194_ _05523_ _00617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06968__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10145_ _04610_ memory\[44\]\[17\] _04944_ _04952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_89_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07383__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10076_ _04915_ _00107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14953_ _01992_ clknet_leaf_35_clk_i memory\[37\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12210__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13904_ _00943_ clknet_leaf_122_clk_i memory\[11\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_85_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14884_ _01923_ clknet_leaf_400_clk_i memory\[35\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07182__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13835_ _00874_ clknet_leaf_205_clk_i memory\[13\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12418__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13766_ _00805_ clknet_leaf_217_clk_i memory\[14\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07145__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10978_ _05024_ memory\[56\]\[9\] _05399_ _05409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_100_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_114_Left_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09834__A2 _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09103__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15505_ _00464_ clknet_leaf_154_clk_i memory\[54\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12717_ memory\[6\]\[17\] memory\[7\]\[17\] _06431_ _02118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08893__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13697_ _03079_ _00766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_80_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15436_ _00395_ clknet_leaf_289_clk_i memory\[52\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08942__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12648_ _03118_ _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_182_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_382_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15367_ _00326_ clknet_leaf_293_clk_i memory\[50\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12579_ memory\[0\]\[15\] memory\[1\]\[15\] memory\[2\]\[15\] memory\[3\]\[15\] _06709_
+ _06779_ _06780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_25_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09837__I _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14318_ _01357_ clknet_leaf_195_clk_i memory\[17\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15298_ _00257_ clknet_leaf_314_clk_i memory\[48\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_41_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14249_ _01288_ clknet_leaf_200_clk_i memory\[15\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_141_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_123_Left_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08810_ _04222_ memory\[25\]\[19\] _04204_ _04223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10712__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09790_ _04763_ _02053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08741_ _03810_ memory\[24\]\[28\] _04168_ _04177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_183_Right_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08672_ _04140_ _01558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12409__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07623_ _03566_ _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_5_Right_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_132_Left_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07554_ _03529_ _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07136__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07485_ _03492_ _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08884__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11342__I _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09224_ _04216_ memory\[31\]\[16\] _04441_ _04448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_157_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10691__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09948__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_180_clk_i clknet_5_29__leaf_clk_i clknet_leaf_180_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_20_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09155_ _04411_ _01770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12374__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07439__I1 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_118_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08106_ _03839_ _01293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_82_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07468__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10443__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_127_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09086_ _04214_ memory\[2\]\[15\] _04369_ _04375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_135_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_141_Left_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08037_ _03798_ memory\[12\]\[22\] _03794_ _03799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_195_clk_i clknet_5_31__leaf_clk_i clknet_leaf_195_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_183_3904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09683__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09061__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12896__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12991__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08299__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09988_ _04589_ memory\[42\]\[7\] _04861_ _04869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08939_ _04285_ _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13696__I0 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Right_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11517__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11950_ memory\[6\]\[6\] memory\[7\]\[6\] _05706_ _06160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07375__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_150_Left_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07931__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10901_ _05368_ _00479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_133_clk_i clknet_5_22__leaf_clk_i clknet_leaf_133_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_28_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11881_ _05710_ _06091_ _06092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_168_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13620_ _05748_ _03003_ _03005_ _03007_ _03008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10832_ _05331_ _00447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13551_ memory\[20\]\[29\] memory\[21\]\[29\] _02368_ _02940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10763_ _05014_ memory\[53\]\[4\] _05290_ _05295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10069__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12820__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11252__I _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_148_clk_i clknet_5_19__leaf_clk_i clknet_leaf_148_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12502_ memory\[4\]\[14\] memory\[5\]\[14\] _06156_ _06704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13482_ _02871_ _02872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_192_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10694_ _05258_ _00382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15221_ _00180_ clknet_leaf_8_clk_i memory\[45\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12433_ memory\[48\]\[13\] memory\[49\]\[13\] memory\[50\]\[13\] memory\[51\]\[13\]
+ _06010_ _06150_ _06636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_30_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15152_ _00111_ clknet_leaf_9_clk_i memory\[43\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12364_ _06149_ _06567_ _06568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14103_ _01142_ clknet_leaf_151_clk_i memory\[63\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11315_ memory\[61\]\[7\] _03146_ _05580_ _05588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15083_ _00042_ clknet_leaf_34_clk_i memory\[41\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12295_ memory\[52\]\[11\] memory\[53\]\[11\] _06143_ _06500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14034_ _01073_ clknet_leaf_139_clk_i memory\[0\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11246_ _03323_ memory\[60\]\[7\] _05543_ _05551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11628__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10532__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11177_ _05514_ _00609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_329_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10128_ _04593_ memory\[44\]\[9\] _04933_ _04943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_141_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10059_ _04906_ _00099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14936_ _01975_ clknet_leaf_71_clk_i memory\[36\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12734__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08937__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_171_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12459__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14867_ _01906_ clknet_leaf_75_clk_i memory\[34\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11363__S _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13818_ _00857_ clknet_leaf_28_clk_i memory\[16\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13064__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12498__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14798_ _01837_ clknet_leaf_50_clk_i memory\[32\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13749_ _03106_ _00791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_139_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07270_ _03374_ _00922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09768__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15419_ _00378_ clknet_leaf_378_clk_i memory\[51\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12194__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07288__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_25__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12922__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09911_ _04828_ _00029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09043__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_130_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09842_ _04579_ memory\[40\]\[2\] _04789_ _04792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11550__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09008__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09773_ _04754_ _02045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06985_ _03194_ memory\[14\]\[22\] _03188_ _03195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_clk_i clknet_5_18__leaf_clk_i clknet_leaf_50_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08724_ _04145_ _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_179_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08847__S _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08655_ _04131_ _01550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12369__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10900__I1 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_53_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07606_ _03557_ _01075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08586_ _04094_ _01518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07109__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_65_clk_i clknet_5_16__leaf_clk_i clknet_leaf_65_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07537_ _03520_ _01043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08857__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07468_ memory\[49\]\[25\] _03361_ _03477_ _03483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09207_ _04199_ memory\[31\]\[8\] _04430_ _04439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07399_ _03444_ _00981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07198__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10416__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09138_ _04402_ _01762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_278_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09282__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09069_ _04197_ memory\[2\]\[7\] _04358_ _04366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_163_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11100_ _03313_ memory\[58\]\[2\] _05471_ _05474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12869__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12080_ _06146_ _06286_ _06287_ _06288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_130_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11031_ _05437_ _00540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12631__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10352__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10344__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output61_I net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_330_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_18_clk_i clknet_5_16__leaf_clk_i clknet_leaf_18_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_189_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10151__I _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15770_ _00729_ clknet_leaf_389_clk_i memory\[62\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12982_ _02358_ _02366_ _02379_ _02380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_51_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07348__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07661__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12787__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14721_ _01760_ clknet_leaf_414_clk_i memory\[30\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11933_ _05677_ _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_19_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14652_ _01691_ clknet_leaf_389_clk_i memory\[28\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13046__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11864_ memory\[56\]\[5\] memory\[57\]\[5\] memory\[58\]\[5\] memory\[59\]\[5\] _05670_
+ _05671_ _06075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_156_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13603_ memory\[40\]\[30\] memory\[41\]\[30\] memory\[42\]\[30\] memory\[43\]\[30\]
+ _05692_ _05694_ _02991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10815_ _05066_ memory\[53\]\[29\] _05312_ _05322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14583_ _01622_ clknet_leaf_79_clk_i memory\[25\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11795_ _06006_ _06007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09588__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13534_ _02344_ _02922_ _02923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08492__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10746_ _05285_ _00407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_11_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13465_ _02319_ _02847_ _02854_ _02855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_11_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10677_ memory\[51\]\[28\] _03211_ _05240_ _05249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_97_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15204_ _00163_ clknet_leaf_399_clk_i memory\[45\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12416_ _06484_ _06619_ _06620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_125_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07028__A2 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09273__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13396_ _02786_ _02787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12652__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11080__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15135_ _00094_ clknet_leaf_439_clk_i memory\[43\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12347_ _06467_ _06544_ _06551_ _06552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__10326__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11780__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07836__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11866__B _06074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15066_ _00025_ clknet_leaf_443_clk_i memory\[40\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12278_ _05759_ _06484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_14017_ _01056_ clknet_leaf_339_clk_i memory\[0\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10262__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11229_ _05541_ _00634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_71_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_71_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08667__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07571__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_37_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12189__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14919_ _01958_ clknet_leaf_20_clk_i memory\[36\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08440_ _04017_ _01449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13037__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_19_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08371_ _03781_ memory\[1\]\[14\] _03976_ _03981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13132__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11599__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07322_ memory\[11\]\[22\] _03355_ _03401_ _03404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09498__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_156_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06915__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07253_ _03205_ _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_171_3660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10437__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_115_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_30_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07184_ _03316_ _00894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_132_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13748__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11771__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07746__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09016__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10172__S _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07578__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09825_ _04781_ _02070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13483__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10900__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09756_ _04744_ _02038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08577__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06968_ _03181_ memory\[14\]\[18\] _03157_ _03182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13276__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08707_ _04159_ _01574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_178_3803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09687_ _04631_ memory\[37\]\[27\] _04700_ _04708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06899_ _03129_ memory\[14\]\[1\] _03126_ _03130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08638_ memory\[23\]\[11\] _03332_ _04121_ _04123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10885__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07750__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08569_ _03775_ memory\[22\]\[11\] _04084_ _04086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10600_ _05056_ memory\[50\]\[24\] _05203_ _05208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11580_ _05693_ _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_119_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12882__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09201__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10531_ _05171_ _00306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13250_ _02167_ _02642_ _05756_ _02643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_88_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09255__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10462_ _05054_ memory\[48\]\[23\] _05131_ _05135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12201_ _05767_ _06400_ _06407_ _06408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_122_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13181_ _02530_ _02545_ _02560_ _02575_ _02576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_10393_ _05098_ _00241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12132_ memory\[22\]\[8\] memory\[23\]\[8\] _06062_ _06340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_92_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11178__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12063_ _06271_ _00738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_53_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07569__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11514__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09871__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11365__I1 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11014_ _05060_ memory\[56\]\[26\] _05421_ _05428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11906__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15822_ _00781_ clknet_leaf_215_clk_i memory\[9\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13267__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15753_ _00712_ clknet_leaf_226_clk_i memory\[62\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12965_ _05669_ _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_73_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13406__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14704_ _01743_ clknet_leaf_89_clk_i memory\[2\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11916_ _05788_ _06126_ _05792_ _06127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15684_ _00643_ clknet_leaf_306_clk_i memory\[60\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12896_ _06480_ _02294_ _06482_ _02295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_158_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13114__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14635_ _01674_ clknet_leaf_185_clk_i memory\[27\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11847_ _05914_ _06054_ _06056_ _06058_ _06059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_129_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12737__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11641__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_136_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14566_ _01605_ clknet_leaf_179_clk_i memory\[25\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11778_ _05788_ _05990_ _05792_ _05991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_144_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09111__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13517_ _05752_ _02905_ _05791_ _02906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10729_ _05047_ memory\[52\]\[20\] _05276_ _05277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14497_ _01536_ clknet_leaf_351_clk_i memory\[23\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11440__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13448_ _05724_ _02837_ _02838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08950__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11053__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09797__I1 _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13379_ _02163_ _02765_ _02767_ _02769_ _02770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_73_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15118_ _00077_ clknet_leaf_21_clk_i memory\[42\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11088__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07940_ _03191_ memory\[19\]\[21\] _03733_ _03735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12271__I _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15049_ _00008_ clknet_leaf_25_clk_i memory\[40\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07871_ _03698_ _01199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11600__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09610_ _04667_ _01969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10720__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_226_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09541_ _04627_ memory\[35\]\[25\] _04617_ _04628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_108_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10867__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09472_ _03134_ _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_188_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08423_ _04008_ _01441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_173_3711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_175_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08354_ _03764_ memory\[1\]\[6\] _03965_ _03972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13430__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09485__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07305_ memory\[11\]\[14\] _03338_ _03390_ _03395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11292__I0 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08285_ _03935_ _01376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09956__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_15_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07236_ memory\[39\]\[20\] _03350_ _03351_ _03352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09237__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12616__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11044__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07167_ _03110_ _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07799__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11744__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07476__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07412__A2 _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07098_ _03226_ _03264_ _03265_ _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_160_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07275__I _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11347__I1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09691__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_31_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09808_ _04772_ _02062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09490__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09739_ _04735_ _02030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_2_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13344__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11525__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10858__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12750_ _06610_ _02150_ _02151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_97_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07723__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11701_ _05655_ _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_16_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12681_ _02082_ _02083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12557__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14420_ _01459_ clknet_leaf_92_clk_i memory\[20\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11632_ _05748_ _05842_ _05844_ _05846_ _05847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_181_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13421__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_428_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09476__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08834__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14351_ _01390_ clknet_leaf_191_clk_i memory\[18\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11563_ _03747_ _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10077__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13302_ _02371_ _02694_ _02373_ _02695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_64_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_94_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10514_ _05162_ _00298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14282_ _01321_ clknet_leaf_182_clk_i memory\[29\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09228__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08770__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11494_ _05667_ _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_126_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13388__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13233_ memory\[24\]\[24\] memory\[25\]\[24\] memory\[26\]\[24\] memory\[27\]\[24\]
+ _02363_ _02502_ _02627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10445_ _05037_ memory\[48\]\[15\] _05120_ _05126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10805__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_175_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11735__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07386__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13164_ _02209_ _02554_ _02556_ _02558_ _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_143_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10376_ _05089_ _00233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11830__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12115_ memory\[46\]\[8\] memory\[47\]\[8\] _05907_ _06323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13095_ _02216_ _02490_ _02491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07185__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11338__I1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12046_ memory\[28\]\[7\] memory\[29\]\[7\] _05915_ _06255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12160__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11636__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10540__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15805_ _00764_ clknet_leaf_287_clk_i memory\[9\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13997_ _01036_ clknet_leaf_228_clk_i memory\[59\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11435__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15736_ _00695_ clknet_leaf_383_clk_i memory\[61\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12948_ memory\[32\]\[20\] memory\[33\]\[20\] memory\[34\]\[20\] memory\[35\]\[20\]
+ _02205_ _02345_ _02346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__13660__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_66_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12467__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15667_ _00626_ clknet_leaf_144_clk_i memory\[5\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_66_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12879_ _02277_ _02278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_103_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11371__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_4033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14618_ _01657_ clknet_leaf_4_clk_i memory\[26\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09467__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15598_ _00557_ clknet_leaf_245_clk_i memory\[57\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11274__I0 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12266__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14549_ _01588_ clknet_leaf_81_clk_i memory\[24\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09776__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08070_ _03754_ memory\[15\]\[1\] _03819_ _03821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_11_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07021_ _03221_ memory\[14\]\[31\] _03125_ _03222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11726__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11821__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12930__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08972_ _04314_ _01684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13479__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07923_ _03166_ memory\[19\]\[13\] _03722_ _03726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_166_3581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07854_ _03689_ _01191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_377_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09016__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07785_ _03163_ memory\[6\]\[12\] _03650_ _03653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09524_ _03186_ _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_17_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08855__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09455_ _04243_ memory\[34\]\[29\] _04560_ _04570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08406_ _03816_ memory\[1\]\[31\] _03964_ _03999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09386_ _04533_ _01879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08337_ _03962_ _01401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11265__I0 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_948 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08130__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08590__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08268_ _03814_ memory\[17\]\[30\] _03892_ _03926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07219_ _03171_ _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_116_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10625__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12904__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08199_ _03889_ _01336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Left_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11717__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10230_ _04627_ memory\[45\]\[25\] _04991_ _04997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06902__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_3946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_186_3957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_424_clk_i clknet_5_0__leaf_clk_i clknet_leaf_424_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10161_ _04960_ _00147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_7_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10092_ _04625_ memory\[43\]\[24\] _04919_ _04924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10360__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13920_ _00959_ clknet_leaf_300_clk_i memory\[8\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07944__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07733__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_439_clk_i clknet_5_0__leaf_clk_i clknet_leaf_439_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13851_ _00890_ clknet_leaf_30_clk_i memory\[13\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_27_Left_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_57_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12802_ _02201_ _02202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13782_ _00821_ clknet_leaf_136_clk_i memory\[14\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_48_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10994_ _05417_ _00523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_48_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15521_ _00480_ clknet_leaf_333_clk_i memory\[55\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12733_ _06450_ _02133_ _06866_ _02134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11191__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15452_ _00411_ clknet_leaf_332_clk_i memory\[53\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12664_ _06863_ _06864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09449__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13245__I1 net56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14403_ _01442_ clknet_leaf_356_clk_i memory\[20\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11615_ memory\[8\]\[1\] memory\[9\]\[1\] memory\[10\]\[1\] memory\[11\]\[1\] _05725_
+ _05726_ _05830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_143_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15383_ _00342_ clknet_leaf_382_clk_i memory\[50\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12595_ _06453_ _06795_ _06796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_53_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09596__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14334_ _01373_ clknet_leaf_350_clk_i memory\[18\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11546_ _05693_ _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_108_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_36_Left_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11008__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14265_ _01304_ clknet_leaf_138_clk_i memory\[15\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11477_ _03116_ _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_150_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13216_ memory\[38\]\[24\] memory\[39\]\[24\] _05662_ _02610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10428_ _05020_ memory\[48\]\[7\] _05109_ _05117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14196_ _01235_ clknet_leaf_104_clk_i memory\[19\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_164_Right_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09621__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12381__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13147_ memory\[8\]\[23\] memory\[9\]\[23\] memory\[10\]\[23\] memory\[11\]\[23\]
+ _02473_ _06721_ _02542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12920__A3 _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10359_ _05080_ _00225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07844__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13078_ memory\[8\]\[22\] memory\[9\]\[22\] memory\[10\]\[22\] memory\[11\]\[22\]
+ _02473_ _06721_ _02474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08188__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12133__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12029_ _06024_ _06233_ _06235_ _06237_ _06238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_174_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_144_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07935__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_68_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_68_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07570_ _03538_ _01058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08675__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15719_ _00678_ clknet_leaf_235_clk_i memory\[61\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_119_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08360__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09240_ _04456_ _01810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09171_ _04231_ memory\[30\]\[23\] _04416_ _04420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12925__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08112__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13492__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08122_ _03806_ memory\[15\]\[26\] _03841_ _03848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_12_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__06923__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__I1 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08053_ _03809_ _01270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10445__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07004_ _03208_ _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_98_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_131_Right_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12372__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10244__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_110_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_164_3529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07754__S _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08955_ _04305_ _01676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_181_3854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11276__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07906_ _03141_ memory\[19\]\[5\] _03711_ _03717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_181_3865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10180__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08886_ _04218_ memory\[26\]\[17\] _04261_ _04269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input23_I data_i[24] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07837_ _03680_ _01183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_123_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08585__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07768_ _03138_ memory\[6\]\[4\] _03639_ _03644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09679__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09507_ _04604_ memory\[35\]\[14\] _04596_ _04605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07699_ _03607_ _01118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09438_ _04561_ _01903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11238__I0 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09369_ _04224_ memory\[33\]\[20\] _04524_ _04525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08103__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11938__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11400_ _03340_ memory\[62\]\[15\] _05627_ _05633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07929__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12380_ _06031_ _06583_ _06584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11959__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08654__I1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11331_ _05596_ _00681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14050_ _01089_ clknet_leaf_303_clk_i memory\[10\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11262_ _05559_ _00649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_363_clk_i clknet_5_9__leaf_clk_i clknet_leaf_363_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_48_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13001_ _02302_ _02390_ _02397_ _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_10213_ _04610_ memory\[45\]\[17\] _04980_ _04988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11193_ _03338_ memory\[5\]\[14\] _05518_ _05523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07090__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_89_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10144_ _04951_ _00139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_89_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_378_clk_i clknet_5_6__leaf_clk_i clknet_leaf_378_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10090__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10075_ _04608_ memory\[43\]\[16\] _04908_ _04915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14952_ _01991_ clknet_leaf_36_clk_i memory\[37\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12210__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07917__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13903_ _00942_ clknet_leaf_202_clk_i memory\[11\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14883_ _01922_ clknet_leaf_428_clk_i memory\[35\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08590__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13834_ _00873_ clknet_leaf_202_clk_i memory\[13\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_5_5__f_clk_i clknet_2_0_0_clk_i clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_301_clk_i clknet_5_14__leaf_clk_i clknet_leaf_301_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xmax_cap72 _03565_ net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_35_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13765_ _00804_ clknet_leaf_275_clk_i memory\[14\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10977_ _05408_ _00515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12809__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08342__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_63_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15504_ _00463_ clknet_leaf_154_clk_i memory\[54\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08294__I _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12716_ _02116_ _02117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13696_ _03315_ memory\[9\]\[3\] _03075_ _03079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12647_ _06846_ _06847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_316_clk_i clknet_5_11__leaf_clk_i clknet_leaf_316_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15435_ _00394_ clknet_leaf_296_clk_i memory\[52\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10329__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12745__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15366_ _00325_ clknet_leaf_293_clk_i memory\[50\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12578_ _03116_ _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09842__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12441__I2 memory\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_15__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14317_ _01356_ clknet_leaf_194_clk_i memory\[17\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11529_ _05741_ _05744_ _05745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10265__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15297_ _00256_ clknet_leaf_329_clk_i memory\[48\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14248_ _01287_ clknet_leaf_200_clk_i memory\[15\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14179_ _01218_ clknet_leaf_341_clk_i memory\[19\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_68_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11096__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08740_ _04176_ _01590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07908__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08671_ memory\[23\]\[27\] _03365_ _04132_ _04140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08581__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11960__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07622_ _03115_ net72 _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__13606__A1 _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07553_ _03227_ _03528_ _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_49_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07484_ _03491_ _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_76_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09223_ _04447_ _01802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06895__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12655__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_20_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09154_ _04214_ memory\[30\]\[15\] _04405_ _04411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08636__I1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08105_ _03789_ memory\[15\]\[18\] _03830_ _03839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12593__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09085_ _04374_ _01737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09964__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08036_ _03193_ _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_141_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11779__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12390__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07072__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09987_ _04868_ _00065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08938_ _04296_ _01668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_93_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08869_ _04201_ memory\[26\]\[9\] _04250_ _04260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_99_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_274_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10900_ memory\[55\]\[4\] _03137_ _05363_ _05368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11880_ memory\[0\]\[5\] memory\[1\]\[5\] memory\[2\]\[5\] memory\[3\]\[5\] _06020_
+ _06090_ _06091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_28_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10831_ _05014_ memory\[54\]\[4\] _05326_ _05331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08324__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11533__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13550_ _02494_ _02934_ _02936_ _02938_ _02939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10762_ _05294_ _00414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10131__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Right_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_137_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12501_ _06411_ _06694_ _06702_ _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_48_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13481_ memory\[28\]\[28\] memory\[29\]\[28\] _02495_ _02871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10693_ _05012_ memory\[52\]\[3\] _05254_ _05258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15220_ _00179_ clknet_leaf_15_clk_i memory\[45\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07659__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12432_ _06146_ _06634_ _06287_ _06635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_180_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__I1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15151_ _00110_ clknet_leaf_19_clk_i memory\[43\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12363_ memory\[48\]\[12\] memory\[49\]\[12\] memory\[50\]\[12\] memory\[51\]\[12\]
+ _06010_ _06150_ _06567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_14102_ _01141_ clknet_leaf_143_clk_i memory\[63\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_22_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11314_ _05587_ _00673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15082_ _00041_ clknet_leaf_33_clk_i memory\[41\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12294_ _06272_ _06494_ _06496_ _06498_ _06499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_105_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12336__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14033_ _01072_ clknet_leaf_109_clk_i memory\[0\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11245_ _05550_ _00641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_20_Right_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10813__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07394__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_56_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11176_ _03321_ memory\[5\]\[6\] _05507_ _05514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11708__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12313__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10127_ _04942_ _00131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10058_ _04591_ memory\[43\]\[8\] _04897_ _04906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14935_ _01974_ clknet_leaf_12_clk_i memory\[36\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_240_clk_i clknet_5_15__leaf_clk_i clknet_leaf_240_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_187_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14866_ _01905_ clknet_leaf_75_clk_i memory\[34\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_72_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13817_ _00856_ clknet_leaf_108_clk_i memory\[16\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11443__I _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14797_ _01836_ clknet_leaf_51_clk_i memory\[32\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12498__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13748_ _03367_ memory\[9\]\[28\] _03097_ _03106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10122__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_255_clk_i clknet_5_24__leaf_clk_i clknet_leaf_255_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_139_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10673__I1 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13679_ memory\[22\]\[31\] memory\[23\]\[31\] _05754_ _03066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13447__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07569__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_wire73_I _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_14_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15418_ _00377_ clknet_leaf_379_clk_i memory\[51\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11599__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_143_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12274__I _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15349_ _00308_ clknet_leaf_150_clk_i memory\[4\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_130_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09784__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_106_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09910_ _04579_ memory\[41\]\[2\] _04825_ _04828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09583__I _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_130_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09841_ _04791_ _02076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10889__A1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09772_ memory\[3\]\[2\] _03131_ _04751_ _04754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06984_ _03193_ _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08723_ _04167_ _01582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_208_clk_i clknet_5_31__leaf_clk_i clknet_leaf_208_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_179_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08554__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11554__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08654_ memory\[23\]\[19\] _03348_ _04121_ _04131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09024__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07605_ _03200_ memory\[0\]\[24\] _03552_ _03557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13054__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_159_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08585_ _03791_ memory\[22\]\[19\] _04084_ _04094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07536_ memory\[59\]\[24\] _03359_ _03515_ _03520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_76_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08863__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12385__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07467_ _03482_ _01011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09206_ _04438_ _01794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07398_ _03206_ memory\[8\]\[26\] _03437_ _03444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09137_ _04197_ memory\[30\]\[7\] _04394_ _04402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09068_ _04365_ _01729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08019_ _03786_ _01259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10633__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09493__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11030_ _05008_ memory\[57\]\[1\] _05435_ _05437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06910__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08103__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12133__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_34_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output54_I net54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07942__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12981_ _02367_ _02370_ _02374_ _02378_ _02379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_51_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_5_23__f_clk_i clknet_2_2_0_clk_i clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_51_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14720_ _01759_ clknet_leaf_418_clk_i memory\[30\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11932_ _05675_ _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08837__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10352__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11863_ _05660_ _06073_ _06001_ _06074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14651_ _01690_ clknet_leaf_4_clk_i memory\[27\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13602_ _05682_ _02989_ _05722_ _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09869__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10814_ _05321_ _00439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10104__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14582_ _01621_ clknet_leaf_84_clk_i memory\[25\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08773__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11794_ memory\[52\]\[4\] memory\[53\]\[4\] _05678_ _06006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10745_ _05064_ memory\[52\]\[28\] _05276_ _05285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12295__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13533_ memory\[32\]\[29\] memory\[33\]\[29\] memory\[34\]\[29\] memory\[35\]\[29\]
+ _05670_ _02345_ _02922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_153_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13429__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13464_ _05768_ _02849_ _02851_ _02853_ _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_11_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10676_ _05248_ _00374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_11_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12415_ memory\[16\]\[12\] memory\[17\]\[12\] memory\[18\]\[12\] memory\[19\]\[12\]
+ _06342_ _06485_ _06619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_15203_ _00162_ clknet_leaf_429_clk_i memory\[45\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11604__I0 memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12094__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13395_ memory\[12\]\[27\] memory\[13\]\[27\] _05769_ _02786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12652__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07188__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12346_ _06476_ _06546_ _06548_ _06550_ _06551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15134_ _00093_ clknet_leaf_440_clk_i memory\[43\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_58_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12309__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_75_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15065_ _00024_ clknet_leaf_3_clk_i memory\[40\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12277_ _06480_ _06481_ _06482_ _06483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_75_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07916__I _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09109__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14016_ _01055_ clknet_leaf_341_clk_i memory\[0\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07036__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11228_ _03373_ memory\[5\]\[31\] _05506_ _05541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13139__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11438__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_71_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11159_ _05504_ _00601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08948__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12168__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08536__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14918_ _01957_ clknet_leaf_35_clk_i memory\[36\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_188_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10894__I1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14849_ _01888_ clknet_leaf_426_clk_i memory\[34\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_194_clk_i clknet_5_31__leaf_clk_i clknet_leaf_194_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08370_ _03980_ _01416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08683__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07321_ _03403_ _00944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12796__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13602__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10646__I1 _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10718__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_154_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12260__A3 _06465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07511__I1 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07299__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07252_ _03362_ _00916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_3661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_222_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_115_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07183_ memory\[39\]\[3\] _03315_ _03309_ _03316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_132_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06931__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_132_clk_i clknet_5_28__leaf_clk_i clknet_leaf_132_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_42_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10453__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12720__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10252__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09824_ memory\[3\]\[27\] _03208_ _04773_ _04781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_147_clk_i clknet_5_22__leaf_clk_i clknet_leaf_147_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07762__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06967_ _03180_ _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09755_ _04631_ memory\[38\]\[27\] _04736_ _04744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11284__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08706_ _03775_ memory\[24\]\[11\] _04157_ _04159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09686_ _04707_ _02005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06898_ _03128_ _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08637_ _04122_ _01541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13659__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08568_ _04085_ _01509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12787__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07519_ memory\[59\]\[16\] _03342_ _03504_ _03511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10637__I1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08499_ _03772_ memory\[21\]\[10\] _04048_ _04049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13004__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07502__I1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12882__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10530_ _05054_ memory\[4\]\[23\] _05167_ _05171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12539__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10461_ _05134_ _00273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12843__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12200_ _05783_ _06402_ _06404_ _06406_ _06407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_44_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13180_ _02358_ _02567_ _02574_ _02575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_126_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10392_ _05052_ memory\[47\]\[22\] _05095_ _05098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12131_ _06338_ _06339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_62_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_36_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12062_ _06270_ net69 _05802_ _06271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_424_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11013_ _05427_ _00532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10573__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07672__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15821_ _00780_ clknet_leaf_214_clk_i memory\[9\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15752_ _00711_ clknet_leaf_225_clk_i memory\[62\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12964_ _06607_ _02361_ _02086_ _02362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09191__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_171_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14703_ _01742_ clknet_leaf_168_clk_i memory\[2\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12570__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11915_ memory\[22\]\[5\] memory\[23\]\[5\] _06062_ _06126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15683_ _00642_ clknet_leaf_322_clk_i memory\[60\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12895_ memory\[22\]\[19\] memory\[23\]\[19\] _06751_ _02294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11922__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14634_ _01673_ clknet_leaf_186_clk_i memory\[27\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11846_ _05921_ _06057_ _06058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_184_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_136_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12322__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11777_ memory\[22\]\[3\] memory\[23\]\[3\] _05789_ _05990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14565_ _01604_ clknet_leaf_408_clk_i memory\[25\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12817__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10538__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13516_ memory\[6\]\[29\] memory\[7\]\[29\] _02322_ _02905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11450__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10728_ _05253_ _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_67_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14496_ _01535_ clknet_leaf_350_clk_i memory\[23\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13447_ memory\[48\]\[28\] memory\[49\]\[28\] memory\[50\]\[28\] memory\[51\]\[28\]
+ _05725_ _05726_ _02837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10659_ _05239_ _00366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13378_ _02170_ _02768_ _02769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__11369__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15117_ _00076_ clknet_leaf_24_clk_i memory\[42\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12329_ memory\[40\]\[11\] memory\[41\]\[11\] memory\[42\]\[11\] memory\[43\]\[11\]
+ _06186_ _06326_ _06534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_110_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_96_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07009__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15048_ _00007_ clknet_leaf_29_clk_i memory\[40\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_64_clk_i clknet_5_16__leaf_clk_i clknet_leaf_64_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_76_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13584__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13750__I0 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07870_ _03187_ memory\[7\]\[20\] _03697_ _03698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10564__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07582__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08509__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_79_clk_i clknet_5_17__leaf_clk_i clknet_leaf_79_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09540_ _03202_ _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_108_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08477__I _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08134__A1 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09471_ _04580_ _01917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08422_ _03764_ memory\[20\]\[6\] _04001_ _04008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_148_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_173_3712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12769__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10619__I1 _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08353_ _03971_ _01408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07304_ _03394_ _00936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_178_Right_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08284_ _03762_ memory\[18\]\[5\] _03929_ _03935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_62_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_11_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_373_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17_clk_i clknet_5_5__leaf_clk_i clknet_leaf_17_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07235_ _03308_ _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12663__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12616__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13194__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07166_ _03302_ _00890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07097_ _03120_ _03122_ _03265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_100_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08588__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07492__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09807_ memory\[3\]\[19\] _03183_ _04762_ _04772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07999_ _03751_ _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11806__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09738_ _04614_ memory\[38\]\[19\] _04725_ _04735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09173__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12552__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09669_ _04698_ _01997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11700_ _05675_ _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_12680_ memory\[28\]\[16\] memory\[29\]\[16\] _06604_ _02082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09212__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11631_ _05760_ _05845_ _05846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10358__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11541__I _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14350_ _01389_ clknet_leaf_196_clk_i memory\[18\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_145_Right_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11562_ _05669_ _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_119_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13301_ memory\[22\]\[25\] memory\[23\]\[25\] _05754_ _02694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10513_ _05037_ memory\[4\]\[15\] _05156_ _05162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14281_ _01320_ clknet_leaf_175_clk_i memory\[29\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_94_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11493_ _05705_ _05707_ _05708_ _05709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_94_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13232_ _02498_ _02625_ _02086_ _02626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_134_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08850__I _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10444_ _05125_ _00265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_118_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11735__A2 _05947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08987__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11189__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13163_ _02216_ _02557_ _02558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10375_ _05035_ memory\[47\]\[14\] _05084_ _05089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10794__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12114_ _05681_ _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09882__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13094_ memory\[40\]\[22\] memory\[41\]\[22\] memory\[42\]\[22\] memory\[43\]\[22\]
+ _06875_ _02217_ _02490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08739__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13732__I0 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12045_ _05731_ _06246_ _06253_ _06254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10546__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12321__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15804_ _00763_ clknet_leaf_283_clk_i memory\[9\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13996_ _01035_ clknet_leaf_227_clk_i memory\[59\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12999__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15735_ _00694_ clknet_leaf_149_clk_i memory\[61\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12947_ _03747_ _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08911__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11652__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11671__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15666_ _00625_ clknet_leaf_141_clk_i memory\[5\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_66_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12878_ memory\[44\]\[19\] memory\[45\]\[19\] _02210_ _02277_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_190_4023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14617_ _01656_ clknet_leaf_79_clk_i memory\[26\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10268__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11829_ _05736_ _06040_ _05739_ _06041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_56_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11451__I _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15597_ _00556_ clknet_leaf_230_clk_i memory\[57\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14548_ _01587_ clknet_leaf_95_clk_i memory\[24\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_112_Right_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13579__S _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12483__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14479_ _01518_ clknet_leaf_175_clk_i memory\[22\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_114_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13176__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07020_ _03220_ _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_102_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08760__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_49_Right_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_149_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08971_ _04235_ memory\[27\]\[25\] _04308_ _04314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13723__I0 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07922_ _03725_ _01223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_166_3571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10731__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07402__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07853_ _03163_ memory\[7\]\[12\] _03686_ _03689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_127_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07784_ _03652_ _01158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_58_Right_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_127_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09523_ _04615_ _01934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_5_4__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09454_ _04569_ _01911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08405_ _03998_ _01433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10178__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09385_ _04241_ memory\[33\]\[28\] _04524_ _04533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08336_ _03814_ memory\[18\]\[30\] _03928_ _03962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08267_ _03925_ _01368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12393__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10906__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_67_Right_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07218_ _03339_ _00905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_41_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08198_ _03812_ memory\[29\]\[29\] _03879_ _03889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08969__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07149_ _03197_ memory\[13\]\[23\] _03290_ _03294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10776__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_186_3958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10160_ _04625_ memory\[44\]\[24\] _04955_ _04960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10091_ _04923_ _00114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10528__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09207__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11536__I _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_76_Right_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13850_ _00889_ clknet_leaf_30_clk_i memory\[13\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_87_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07950__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09146__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12801_ memory\[36\]\[18\] memory\[37\]\[18\] _06447_ _02201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_187_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13781_ _00820_ clknet_leaf_135_clk_i memory\[14\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12568__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10993_ _05039_ memory\[56\]\[16\] _05410_ _05417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_48_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_44_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15520_ _00479_ clknet_leaf_333_clk_i memory\[55\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12732_ memory\[38\]\[17\] memory\[39\]\[17\] _06728_ _02133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15451_ _00410_ clknet_leaf_374_clk_i memory\[52\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10088__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12663_ memory\[36\]\[16\] memory\[37\]\[16\] _06447_ _06863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14402_ _01441_ clknet_leaf_358_clk_i memory\[20\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09877__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11614_ _05719_ _05828_ _05722_ _05829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15382_ _00341_ clknet_5_7__leaf_clk_i memory\[50\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12594_ memory\[32\]\[15\] memory\[33\]\[15\] memory\[34\]\[15\] memory\[35\]\[15\]
+ _06314_ _06454_ _06795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_136_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_85_Right_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14333_ _01372_ clknet_leaf_363_clk_i memory\[18\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11545_ _05691_ _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_25_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07880__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14264_ _01303_ clknet_leaf_140_clk_i memory\[15\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11476_ _05691_ _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA_clkbuf_leaf_269_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10427_ _05116_ _00257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13215_ _02608_ _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_122_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14195_ _01234_ clknet_leaf_102_clk_i memory\[19\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10767__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07632__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13146_ _06717_ _02540_ _02195_ _02541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_21_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10358_ _05018_ memory\[47\]\[6\] _05073_ _05080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13077_ _05669_ _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_100_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10519__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10289_ _03168_ _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_100_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13330__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Right_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09385__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_321_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09117__S _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12028_ _06031_ _06236_ _06237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08021__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11446__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08956__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_68_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09137__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13979_ _01018_ clknet_leaf_379_clk_i memory\[49\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_122_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11644__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15718_ _00677_ clknet_leaf_237_clk_i memory\[61\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15649_ _00608_ clknet_leaf_369_clk_i memory\[5\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09170_ _04419_ _01777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08691__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_1_Left_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08121_ _03847_ _01300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_161_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13492__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13610__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10726__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13149__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08052_ _03808_ memory\[12\]\[27\] _03794_ _03809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07003_ net26 _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_168_3611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12941__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08954_ _04218_ memory\[27\]\[17\] _04297_ _04305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_4_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_181_3855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07905_ _03716_ _01215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_181_3866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08885_ _04268_ _01643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07836_ _03138_ memory\[7\]\[4\] _03675_ _03680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12896__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07770__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_input16_I data_i[18] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07767_ _03643_ _01150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11292__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09506_ _03168_ _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_17_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07698_ _03135_ memory\[63\]\[3\] _03603_ _03607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09437_ _04224_ memory\[34\]\[20\] _04560_ _04561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_23_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09368_ _04501_ _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_152_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08319_ _03953_ _01392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_151_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12060__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09299_ _04487_ _01838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10997__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11330_ memory\[61\]\[14\] _03168_ _05591_ _05596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06913__I net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_270_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11261_ _03338_ memory\[60\]\[14\] _05554_ _05559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10749__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10212_ _04987_ _00171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13000_ _06831_ _02392_ _02394_ _02396_ _02397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_11192_ _05522_ _00616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11975__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10143_ _04608_ memory\[44\]\[16\] _04944_ _04951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10371__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10074_ _04914_ _00106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14951_ _01990_ clknet_leaf_20_clk_i memory\[37\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11174__I0 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13902_ _00941_ clknet_leaf_203_clk_i memory\[11\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11874__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14882_ _01921_ clknet_leaf_429_clk_i memory\[35\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08776__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07680__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09119__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13833_ _00872_ clknet_leaf_215_clk_i memory\[13\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13764_ _00803_ clknet_leaf_276_clk_i memory\[14\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_74_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10976_ _05022_ memory\[56\]\[8\] _05399_ _05408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_63_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15503_ _00462_ clknet_leaf_242_clk_i memory\[54\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12715_ memory\[4\]\[17\] memory\[5\]\[17\] _06845_ _02116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13695_ _03078_ _00765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_80_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13379__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15434_ _00393_ clknet_leaf_297_clk_i memory\[52\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12646_ memory\[4\]\[16\] memory\[5\]\[16\] _06845_ _06846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12051__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15365_ _00324_ clknet_leaf_313_clk_i memory\[50\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10546__S _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12577_ _06159_ _06777_ _06707_ _06778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14316_ _01355_ clknet_leaf_193_clk_i memory\[17\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_740 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07853__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11528_ memory\[32\]\[0\] memory\[33\]\[0\] memory\[34\]\[0\] memory\[35\]\[0\] _05742_
+ _05743_ _05744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_124_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15296_ _00255_ clknet_leaf_329_clk_i memory\[48\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14247_ _01286_ clknet_leaf_218_clk_i memory\[15\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10345__I _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12761__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11459_ _05652_ _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_110_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07855__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_78_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07605__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14178_ _01217_ clknet_leaf_344_clk_i memory\[19\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11377__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10281__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13129_ _02523_ _02524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09358__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I data_i[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13592__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08670_ _04139_ _01557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11865__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07590__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07621_ _03123_ _03375_ _03565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_75_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13605__B _02990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11960__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07552_ _03112_ _03114_ _03528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__11617__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13162__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12001__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07483_ _03376_ _03490_ _03491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_159_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_423_clk_i clknet_5_0__leaf_clk_i clknet_leaf_423_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_158_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09222_ _04214_ memory\[31\]\[15\] _04441_ _04447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_29_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09153_ _04410_ _01769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08097__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10456__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08104_ _03838_ _01292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09084_ _04212_ memory\[2\]\[14\] _04369_ _04374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07844__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_135_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_438_clk_i clknet_5_0__leaf_clk_i clknet_leaf_438_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_135_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08035_ _03797_ _01264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_142_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10255__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12671__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12345__A2 _06549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13542__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11779__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_55_Left_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09986_ _04587_ memory\[42\]\[6\] _04861_ _04868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09980__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08937_ _04201_ memory\[27\]\[9\] _04286_ _04296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10108__A1 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11156__I0 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08021__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11856__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08596__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_217_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08868_ _04259_ _01635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07819_ _03670_ _01175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08799_ _04215_ _01610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_28_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10830_ _05330_ _00446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07005__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_64_Left_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10761_ _05012_ memory\[53\]\[3\] _05290_ _05294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12500_ _06142_ _06696_ _06698_ _06701_ _06702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_192_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10692_ _05257_ _00381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13480_ _02336_ _02862_ _02869_ _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_109_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13250__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12431_ memory\[54\]\[13\] memory\[55\]\[13\] _06421_ _06634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12645__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09824__I1 _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_35_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15150_ _00109_ clknet_leaf_21_clk_i memory\[43\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12362_ _06146_ _06565_ _06287_ _06566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_14101_ _01140_ clknet_leaf_143_clk_i memory\[63\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13677__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11313_ memory\[61\]\[6\] _03143_ _05580_ _05587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15081_ _00040_ clknet_leaf_25_clk_i memory\[41\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12293_ _06279_ _06497_ _06498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_73_Left_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09588__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14032_ _01071_ clknet_leaf_138_clk_i memory\[0\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11244_ _03321_ memory\[60\]\[6\] _05543_ _05550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11197__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_56_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08260__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11175_ _05513_ _00608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09890__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12719__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10126_ _04591_ memory\[44\]\[8\] _04933_ _04942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08012__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13392__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10057_ _04905_ _00098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11847__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14934_ _01973_ clknet_leaf_13_clk_i memory\[36\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_101_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_37_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14865_ _01904_ clknet_leaf_77_clk_i memory\[34\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_82_Left_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13816_ _00855_ clknet_leaf_109_clk_i memory\[16\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14796_ _01835_ clknet_leaf_52_clk_i memory\[32\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13747_ _03105_ _00790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10959_ _05398_ _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_2_3_0_clk_i clknet_0_clk_i clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_139_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11660__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_419_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13678_ _03064_ _03065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_57_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13447__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15417_ _00376_ clknet_leaf_384_clk_i memory\[51\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12629_ _06279_ _06828_ _06829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_14_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15348_ _00307_ clknet_leaf_142_clk_i memory\[4\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_117_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_91_Left_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15279_ _00238_ clknet_leaf_273_clk_i memory\[47\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_166_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13524__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09579__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_113_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_113_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09840_ _04577_ memory\[40\]\[1\] _04789_ _04791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_130_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11630__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10889__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09771_ _04753_ _02044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11138__I0 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06983_ net21 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_20_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11835__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08722_ _03791_ memory\[24\]\[19\] _04157_ _04167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08003__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11838__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09305__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09751__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08653_ _04130_ _01549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13335__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07604_ _03556_ _01074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08584_ _04093_ _01517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_362_clk_i clknet_5_9__leaf_clk_i clknet_leaf_362_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_88_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07535_ _03519_ _01042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_176_3754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11570__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07466_ memory\[49\]\[24\] _03359_ _03477_ _03482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09205_ _04197_ memory\[31\]\[7\] _04430_ _04438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12015__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10186__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07690__A1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07397_ _03443_ _00980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_377_clk_i clknet_5_3__leaf_clk_i clknet_leaf_377_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_162_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09136_ _04401_ _01761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13497__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09067_ _04195_ memory\[2\]\[6\] _04358_ _04365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_load_slew74_I net75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_300_clk_i clknet_5_14__leaf_clk_i clknet_leaf_300_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08018_ _03785_ memory\[12\]\[16\] _03773_ _03786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12414__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11377__I0 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09990__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11129__I0 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_34_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09969_ _04858_ _00057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_315_clk_i clknet_5_10__leaf_clk_i clknet_leaf_315_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11745__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11829__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12980_ _02375_ _02377_ _02378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_368_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output47_I net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_51_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11931_ _05654_ _06135_ _06137_ _06140_ _06141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_169_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11544__I _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14650_ _01689_ clknet_leaf_4_clk_i memory\[27\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11862_ memory\[62\]\[5\] memory\[63\]\[5\] _05868_ _06073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13046__A3 _02442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13601_ memory\[46\]\[30\] memory\[47\]\[30\] _02487_ _02989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_185_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10813_ _05064_ memory\[53\]\[28\] _05312_ _05321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12576__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14581_ _01620_ clknet_leaf_80_clk_i memory\[25\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11688__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11793_ _05654_ _05999_ _06002_ _06004_ _06005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_95_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13532_ _02341_ _02920_ _05708_ _02921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_420_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10744_ _05284_ _00406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13429__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12006__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13463_ _05777_ _02852_ _02853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10096__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10675_ memory\[51\]\[27\] _03208_ _05240_ _05248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15202_ _00161_ clknet_leaf_432_clk_i memory\[45\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_11_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07808__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12414_ _06480_ _06617_ _06482_ _06618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_97_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13394_ _05747_ _02780_ _02782_ _02784_ _02785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_140_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15133_ _00092_ clknet_leaf_434_clk_i memory\[43\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_58_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12345_ _06484_ _06549_ _06550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07284__I1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_26_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15064_ _00023_ clknet_leaf_7_clk_i memory\[40\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12276_ _05791_ _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_142_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14015_ _01054_ clknet_leaf_365_clk_i memory\[0\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08233__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11227_ _05540_ _00633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11158_ _03371_ memory\[58\]\[30\] _05470_ _05504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11655__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10109_ _04932_ _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12168__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11089_ _05467_ _00568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09125__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14917_ _01956_ clknet_leaf_431_clk_i memory\[36\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11454__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_159_Right_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_76_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14848_ _01887_ clknet_leaf_422_clk_i memory\[34\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_19_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_19_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_92_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14779_ _01818_ clknet_leaf_1_clk_i memory\[31\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_193_4076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11390__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07320_ memory\[11\]\[21\] _03353_ _03401_ _03403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08763__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_154_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07251_ memory\[39\]\[25\] _03361_ _03351_ _03362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12285__I _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_171_3662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09795__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07182_ _03134_ _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_115_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_30_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08472__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13110__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_952 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12234__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08224__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09823_ _04780_ _02069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_129_Left_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09754_ _04743_ _02037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06966_ net16 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09035__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13276__A3 _02668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09724__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08705_ _04158_ _01573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09685_ _04629_ memory\[37\]\[26\] _04700_ _04707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06897_ net18 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_126_Right_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_179_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08636_ memory\[23\]\[10\] _03329_ _04121_ _04122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08874__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13659__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12236__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08567_ _03772_ memory\[22\]\[10\] _04084_ _04085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10098__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07518_ _03510_ _01034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08498_ _04036_ _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_138_Left_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_134_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07449_ memory\[49\]\[16\] _03342_ _03466_ _03473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10460_ _05052_ memory\[48\]\[22\] _05131_ _05134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09119_ _04247_ memory\[2\]\[31\] _04357_ _04392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07266__I1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10644__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10391_ _05097_ _00240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_1315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12130_ memory\[20\]\[8\] memory\[21\]\[8\] _05785_ _06338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06921__I net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08114__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12061_ _06224_ _06239_ _06254_ _06269_ _06270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_EDGE_ROW_147_Left_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_53_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10022__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_254_clk_i clknet_5_24__leaf_clk_i clknet_leaf_254_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11012_ _05058_ memory\[56\]\[25\] _05421_ _05427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15820_ _00779_ clknet_leaf_213_clk_i memory\[9\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09715__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15751_ _00710_ clknet_leaf_226_clk_i memory\[62\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12963_ memory\[30\]\[20\] memory\[31\]\[20\] _02084_ _02361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13690__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_269_clk_i clknet_5_13__leaf_clk_i clknet_leaf_269_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_114_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14702_ _01741_ clknet_leaf_169_clk_i memory\[2\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11914_ _06124_ _06125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15682_ _00641_ clknet_leaf_320_clk_i memory\[60\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12570__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12894_ _02292_ _02293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_16_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14633_ _01672_ clknet_leaf_181_clk_i memory\[27\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12227__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_16_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11845_ memory\[24\]\[4\] memory\[25\]\[4\] memory\[26\]\[4\] memory\[27\]\[4\] _05778_
+ _05922_ _06057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10819__S _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_156_Left_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12322__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_28_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14564_ _01603_ clknet_leaf_407_clk_i memory\[25\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11776_ _05988_ _05989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_55_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13515_ _02903_ _02904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10618__I _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10727_ _05275_ _00398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14495_ _01534_ clknet_leaf_351_clk_i memory\[23\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_24_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13446_ _05719_ _02835_ _05739_ _02836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_82_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10658_ memory\[51\]\[19\] _03183_ _05229_ _05239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_207_clk_i clknet_5_31__leaf_clk_i clknet_leaf_207_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_183_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08454__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12833__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10554__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07257__I1 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_495 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13377_ memory\[56\]\[27\] memory\[57\]\[27\] memory\[58\]\[27\] memory\[59\]\[27\]
+ _05711_ _02171_ _02768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_106_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10589_ _05045_ memory\[50\]\[19\] _05192_ _05202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15116_ _00075_ clknet_leaf_2_clk_i memory\[42\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12328_ _06322_ _06532_ _06461_ _06533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08024__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_39_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11449__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08206__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15047_ _00006_ clknet_leaf_22_clk_i memory\[40\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12259_ _06318_ _06459_ _06462_ _06464_ _06465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_43_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10013__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07863__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09954__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11385__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_0_clk_i clk_i clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_78_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12466__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11184__I _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08134__A2 _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09470_ _04579_ memory\[35\]\[2\] _04575_ _04580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08421_ _04007_ _01440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10729__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06940__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08352_ _03762_ memory\[1\]\[5\] _03965_ _03971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13510__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07103__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07303_ memory\[11\]\[13\] _03336_ _03390_ _03394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07496__I1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08283_ _03934_ _01375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08693__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12944__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_316_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07234_ _03186_ _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_143_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08445__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07165_ _03221_ memory\[13\]\[31\] _03267_ _03302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07248__I1 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10464__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07096_ _03117_ _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_4
XFILLER_0_125_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09945__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_31_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09806_ _04771_ _02061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13329__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07420__I1 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07998_ _03155_ _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09737_ _04734_ _02029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06949_ _03167_ _00808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12552__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09668_ _04612_ memory\[37\]\[18\] _04689_ _04698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08619_ memory\[23\]\[2\] _03313_ _04110_ _04113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12209__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06931__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09599_ _04661_ _01964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11630_ memory\[40\]\[1\] memory\[41\]\[1\] memory\[42\]\[1\] memory\[43\]\[1\] _05761_
+ _05762_ _05845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07013__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11561_ _05689_ _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_92_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13300_ _02692_ _02693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_24_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_64_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07948__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10512_ _05161_ _00297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14280_ _01319_ clknet_leaf_182_clk_i memory\[29\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11492_ _05686_ _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_165_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13231_ memory\[30\]\[24\] memory\[31\]\[24\] _02084_ _02625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10443_ _05035_ memory\[48\]\[14\] _05120_ _05125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07239__I1 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13162_ memory\[40\]\[23\] memory\[41\]\[23\] memory\[42\]\[23\] memory\[43\]\[23\]
+ _06875_ _02217_ _02557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_62_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10374_ _05088_ _00232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_40_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_193_clk_i clknet_5_31__leaf_clk_i clknet_leaf_193_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12113_ _06320_ _06321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_27_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13093_ _02213_ _02488_ _02352_ _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08779__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12044_ _05748_ _06248_ _06250_ _06252_ _06253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12696__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09561__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15803_ _00762_ clknet_leaf_26_clk_i net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13995_ _01034_ clknet_leaf_230_clk_i memory\[59\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15734_ _00693_ clknet_leaf_149_clk_i memory\[61\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12946_ _05667_ _02344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__09403__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_88_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_131_clk_i clknet_5_29__leaf_clk_i clknet_leaf_131_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15665_ _00624_ clknet_leaf_144_clk_i memory\[5\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11671__A2 _05884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12877_ _06446_ _02271_ _02273_ _02275_ _02276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_103_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14616_ _01655_ clknet_leaf_77_clk_i memory\[26\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_190_4035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11828_ memory\[38\]\[4\] memory\[39\]\[4\] _06039_ _06040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15596_ _00555_ clknet_leaf_227_clk_i memory\[57\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12049__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14547_ _01586_ clknet_leaf_95_clk_i memory\[24\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07478__I1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11759_ _05732_ _05967_ _05969_ _05971_ _05972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12620__A1 _06774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_146_clk_i clknet_5_22__leaf_clk_i clknet_leaf_146_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10482__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14478_ _01517_ clknet_leaf_197_clk_i memory\[22\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13429_ memory\[16\]\[27\] memory\[17\]\[27\] memory\[18\]\[27\] memory\[19\]\[27\]
+ _02233_ _02376_ _02820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10284__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10234__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06989__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10083__I _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_149_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08970_ _04313_ _01683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_149_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08689__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09927__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07921_ _03163_ memory\[19\]\[12\] _03722_ _03725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12687__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07852_ _03688_ _01190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_127_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput1 address_i[0] net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_07783_ _03160_ memory\[6\]\[11\] _03650_ _03652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11843__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09522_ _04614_ memory\[35\]\[19\] _04596_ _04615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_189_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09313__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13343__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09453_ _04241_ memory\[34\]\[28\] _04560_ _04569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08404_ _03814_ memory\[1\]\[30\] _03964_ _03998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_47_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09384_ _04532_ _01878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08335_ _03961_ _01400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10258__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12611__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07768__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08266_ _03812_ memory\[17\]\[29\] _03915_ _03925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08418__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07217_ memory\[39\]\[14\] _03338_ _03330_ _03339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10194__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08197_ _03888_ _01335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07148_ _03293_ _00881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_186_3948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_186_3959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07079_ _03255_ _00850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09918__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10090_ _04623_ memory\[43\]\[23\] _04919_ _04923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_7_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12678__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11753__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12800_ _06428_ _02190_ _02199_ _02200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_87_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13780_ _00819_ clknet_leaf_113_clk_i memory\[14\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07157__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10992_ _05416_ _00522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_48_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12731_ _02131_ _02132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12648__I _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10369__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11552__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15450_ _00409_ clknet_leaf_270_clk_i memory\[52\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12662_ _06428_ _06854_ _06861_ _06862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_139_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_clk_i clknet_5_16__leaf_clk_i clknet_leaf_63_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14401_ _01440_ clknet_leaf_352_clk_i memory\[20\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11613_ memory\[14\]\[1\] memory\[15\]\[1\] _05720_ _05828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12584__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12602__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15381_ _00340_ clknet_leaf_155_clk_i memory\[50\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12593_ _06450_ _06793_ _06177_ _06794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_108_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07678__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14332_ _01371_ clknet_leaf_363_clk_i memory\[18\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10464__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11544_ _05759_ _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_92_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14263_ _01302_ clknet_leaf_112_clk_i memory\[15\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_78_clk_i clknet_5_17__leaf_clk_i clknet_leaf_78_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11475_ _03119_ _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_21_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13214_ memory\[36\]\[24\] memory\[37\]\[24\] _02338_ _02608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10426_ _05018_ memory\[48\]\[6\] _05109_ _05116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14194_ _01233_ clknet_leaf_102_clk_i memory\[19\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09082__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13145_ memory\[14\]\[23\] memory\[15\]\[23\] _02193_ _02540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10357_ _05079_ _00224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13076_ _06717_ _02471_ _02195_ _02472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13428__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10288_ _05034_ _00200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12027_ memory\[8\]\[7\] memory\[9\]\[7\] memory\[10\]\[7\] memory\[11\]\[7\] _05893_
+ _06032_ _06236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07396__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_16_clk_i clknet_5_5__leaf_clk_i clknet_leaf_16_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_105_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13978_ _01017_ clknet_leaf_380_clk_i memory\[49\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09133__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12929_ _06844_ _02321_ _02324_ _02326_ _02327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15717_ _00676_ clknet_leaf_306_clk_i memory\[61\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11462__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15648_ _00607_ clknet_leaf_369_clk_i memory\[5\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15579_ _00538_ clknet_leaf_374_clk_i memory\[56\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08120_ _03804_ memory\[15\]\[25\] _03841_ _03847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07588__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08051_ _03208_ _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07002_ _03207_ _00821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10207__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09073__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08820__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_122_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08953_ _04304_ _01675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08212__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_110_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07904_ _03138_ memory\[19\]\[4\] _03711_ _03716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08884_ _04216_ memory\[26\]\[16\] _04261_ _04268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_181_3856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_102_Left_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_37_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08011__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07835_ _03679_ _01182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07766_ _03135_ memory\[6\]\[3\] _03639_ _03643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09043__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_8_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09505_ _04603_ _01928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12832__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07697_ _03606_ _01117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09978__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09436_ _04537_ _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08882__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_43_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09367_ _04523_ _01870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_23_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10917__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07498__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08318_ _03796_ memory\[18\]\[21\] _03951_ _03953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09298_ _04222_ memory\[32\]\[19\] _04477_ _04487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_213_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08249_ _03916_ _01359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11260_ _05558_ _00648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10211_ _04608_ memory\[45\]\[16\] _04980_ _04987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_5_17__f_clk_i clknet_2_2_0_clk_i clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_127_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10652__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11191_ _03336_ memory\[5\]\[13\] _05518_ _05522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09218__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10142_ _04950_ _00138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08122__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12152__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10073_ _04606_ memory\[43\]\[15\] _04908_ _04914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14950_ _01989_ clknet_leaf_35_clk_i memory\[37\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13901_ _00940_ clknet_leaf_214_clk_i memory\[11\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14881_ _01920_ clknet_leaf_420_clk_i memory\[35\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10921__I1 _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13832_ _00871_ clknet_leaf_216_clk_i memory\[13\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13076__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08878__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12378__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13763_ _00802_ clknet_leaf_279_clk_i memory\[14\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10975_ _05407_ _00514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_63_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_63_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09888__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15502_ _00461_ clknet_leaf_241_clk_i memory\[54\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12714_ _06411_ _02107_ _02114_ _02115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08792__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13694_ _03313_ memory\[9\]\[2\] _03075_ _03078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15433_ _00392_ clknet_leaf_297_clk_i memory\[52\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12645_ _05701_ _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_80_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10827__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10437__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15364_ _00323_ clknet_leaf_313_clk_i memory\[50\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12576_ memory\[6\]\[15\] memory\[7\]\[15\] _06431_ _06777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07201__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14315_ _01354_ clknet_leaf_194_clk_i memory\[17\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11527_ _03747_ _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_15295_ _00254_ clknet_leaf_347_clk_i memory\[48\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14246_ _01285_ clknet_leaf_218_clk_i memory\[15\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11458_ _05654_ _05658_ _05666_ _05673_ _05674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__09055__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13000__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07000__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_78_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10409_ _05106_ _00249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14177_ _01216_ clknet_leaf_343_clk_i memory\[19\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10562__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11389_ _05615_ _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_21_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13128_ memory\[52\]\[23\] memory\[53\]\[23\] _06832_ _02523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_163_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_415_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13059_ _02454_ _02455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07369__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08967__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12997__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07620_ _03564_ _01082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08766__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_162_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07551_ _03527_ _01050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13162__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08869__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12665__I1 memory\[39\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_9_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07482_ _03113_ _03450_ _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_75_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09221_ _04446_ _01801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10737__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10428__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09152_ _04212_ memory\[30\]\[14\] _04405_ _04410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09294__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07111__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08103_ _03787_ memory\[15\]\[17\] _03830_ _03838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09083_ _04373_ _01736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_140_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08034_ _03796_ memory\[12\]\[21\] _03794_ _03797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_135_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_13_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10472__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_87_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10600__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09985_ _04867_ _00064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Left_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08936_ _04295_ _01667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10108__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07781__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08867_ _04199_ memory\[26\]\[8\] _04250_ _04259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07818_ _03212_ memory\[6\]\[28\] _03661_ _03670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08798_ _04214_ memory\[25\]\[15\] _04204_ _04215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_28_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07749_ _03633_ _01142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_28_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10760_ _05293_ _00413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09501__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09419_ _04551_ _01894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10691_ _05010_ memory\[52\]\[2\] _05254_ _05257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12430_ _06632_ _06633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_63_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09300__I _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07021__S _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_364_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11092__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12361_ memory\[54\]\[12\] memory\[55\]\[12\] _06421_ _06565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14100_ _01139_ clknet_leaf_146_clk_i memory\[63\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11792__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07956__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11312_ _05586_ _00672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09037__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11986__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15080_ _00039_ clknet_leaf_28_clk_i memory\[41\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12292_ memory\[56\]\[11\] memory\[57\]\[11\] memory\[58\]\[11\] memory\[59\]\[11\]
+ _06138_ _06280_ _06497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_14031_ _01070_ clknet_leaf_249_clk_i memory\[0\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11243_ _05549_ _00640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07599__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11174_ _03319_ memory\[5\]\[5\] _05507_ _05513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_56_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10125_ _04941_ _00130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12719__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13297__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_141_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13392__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10056_ _04589_ memory\[43\]\[7\] _04897_ _04905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14933_ _01972_ clknet_leaf_73_clk_i memory\[36\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12102__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14864_ _01903_ clknet_leaf_77_clk_i memory\[34\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13815_ _00854_ clknet_leaf_111_clk_i memory\[16\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14795_ _01834_ clknet_leaf_53_clk_i memory\[32\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13746_ _03365_ memory\[9\]\[27\] _03097_ _03105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10958_ _03227_ _03490_ _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_168_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09411__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_139_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13677_ memory\[20\]\[31\] memory\[21\]\[31\] _05749_ _03064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10889_ _03306_ _03451_ _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_0_183_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12628_ memory\[56\]\[16\] memory\[57\]\[16\] memory\[58\]\[16\] memory\[59\]\[16\]
+ _06827_ _06280_ _06828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15416_ _00375_ clknet_leaf_384_clk_i memory\[51\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08027__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_14_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15347_ _00306_ clknet_leaf_143_clk_i memory\[4\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12559_ memory\[60\]\[15\] memory\[61\]\[15\] _06273_ _06760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11783__A1 _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_152_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15278_ _00237_ clknet_leaf_272_clk_i memory\[47\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_109_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_9_Right_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_112_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14229_ _01268_ clknet_leaf_112_clk_i memory\[12\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_113_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07665__I _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_130_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11630__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_107_Right_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09770_ memory\[3\]\[1\] _03128_ _04751_ _04753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06982_ _03192_ _00816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08697__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08721_ _04166_ _01581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08652_ memory\[23\]\[18\] _03346_ _04121_ _04130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07762__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07603_ _03197_ memory\[0\]\[23\] _03552_ _03556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08583_ _03789_ memory\[22\]\[18\] _04084_ _04093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11851__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07534_ memory\[59\]\[23\] _03357_ _03515_ _03519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_176_3755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__S _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07465_ _03481_ _01010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09204_ _04437_ _01793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13212__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09267__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07396_ _03203_ memory\[8\]\[25\] _03437_ _03443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07690__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11074__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09135_ _04195_ memory\[30\]\[6\] _04394_ _04401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11774__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07776__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09066_ _04364_ _01728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_5_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08017_ _03174_ _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_130_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07575__I _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09968_ _04637_ memory\[41\]\[30\] _04824_ _04858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08919_ _04181_ memory\[27\]\[0\] _04286_ _04287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08400__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09899_ _04821_ _00024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_51_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11930_ _05668_ _06139_ _06140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_51_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_174_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11861_ _06071_ _06072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_13600_ _02987_ _02988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10812_ _05320_ _00438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14580_ _01619_ clknet_leaf_95_clk_i memory\[25\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11792_ _05668_ _06003_ _06004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11688__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11301__I1 _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13531_ memory\[38\]\[29\] memory\[39\]\[29\] _05662_ _02920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10743_ _05062_ memory\[52\]\[27\] _05276_ _05284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10377__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13462_ memory\[8\]\[28\] memory\[9\]\[28\] memory\[10\]\[28\] memory\[11\]\[28\]
+ _02473_ _05779_ _02852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_54_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10674_ _05247_ _00373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_129_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15201_ _00160_ clknet_leaf_423_clk_i memory\[45\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12413_ memory\[22\]\[12\] memory\[23\]\[12\] _06062_ _06617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11065__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13393_ _05759_ _02783_ _02784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12592__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11765__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15132_ _00091_ clknet_leaf_440_clk_i memory\[43\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07686__S _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12344_ memory\[16\]\[11\] memory\[17\]\[11\] memory\[18\]\[11\] memory\[19\]\[11\]
+ _06342_ _06485_ _06549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_110_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_65_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15063_ _00022_ clknet_leaf_9_clk_i memory\[40\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12275_ memory\[22\]\[10\] memory\[23\]\[10\] _06062_ _06481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_75_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13062__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07485__I _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14014_ _01053_ clknet_leaf_365_clk_i memory\[0\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11226_ _03371_ memory\[5\]\[30\] _05506_ _05540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09430__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12190__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_422_clk_i clknet_5_0__leaf_clk_i clknet_leaf_422_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11157_ _05503_ _00600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10108_ _03750_ _04787_ _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_11088_ _05066_ memory\[57\]\[29\] _05457_ _05467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10879__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10039_ _04895_ _00090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14916_ _01955_ clknet_leaf_430_clk_i memory\[36\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07744__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_437_clk_i clknet_5_0__leaf_clk_i clknet_leaf_437_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_188_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14847_ _01886_ clknet_leaf_424_clk_i memory\[34\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_19_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_35_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13442__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14778_ _01817_ clknet_leaf_2_clk_i memory\[31\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_193_4077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09141__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13729_ _03348_ memory\[9\]\[19\] _03086_ _03096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10287__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11470__I _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_154_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_154_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07250_ _03202_ _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_116_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09249__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12628__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07181_ _03314_ _00893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11756__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10803__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_132_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11359__I1 _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12020__I2 memory\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09822_ memory\[3\]\[26\] _03205_ _04773_ _04780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_312_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09753_ _04629_ memory\[38\]\[26\] _04736_ _04743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06965_ _03179_ _00812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08220__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08704_ _03772_ memory\[24\]\[10\] _04157_ _04158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09684_ _04706_ _02004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06896_ _03127_ _00795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08635_ _04109_ _04121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_94_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08566_ _04072_ _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_138_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13433__A1 _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09488__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12867__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__S _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07517_ memory\[59\]\[15\] _03340_ _03504_ _03510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08497_ _04047_ _01476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11995__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09986__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08890__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07448_ _03472_ _01002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_853 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07379_ _03178_ memory\[8\]\[17\] _03426_ _03434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10925__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13301__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09118_ _04391_ _01753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_161_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09660__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10390_ _05050_ memory\[47\]\[21\] _05095_ _05097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12425__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09049_ _04245_ memory\[28\]\[30\] _04321_ _04355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12060_ _05767_ _06261_ _06268_ _06269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_53_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11011_ _05426_ _00531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09226__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08130__S _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12160__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12962_ _02359_ _02360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15750_ _00709_ clknet_leaf_222_clk_i memory\[62\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_5_24__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14701_ _01740_ clknet_leaf_176_clk_i memory\[2\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11913_ memory\[20\]\[5\] memory\[21\]\[5\] _05785_ _06124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_59_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12893_ memory\[20\]\[19\] memory\[21\]\[19\] _06477_ _02292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15681_ _00640_ clknet_leaf_323_clk_i memory\[60\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11491__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14632_ _01671_ clknet_leaf_180_clk_i memory\[27\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11844_ _05918_ _06055_ _05775_ _06056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_16_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13424__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09479__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11286__I0 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14563_ _01602_ clknet_leaf_413_clk_i memory\[25\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_136_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11775_ memory\[20\]\[3\] memory\[21\]\[3\] _05785_ _05988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11986__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09896__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10726_ _05045_ memory\[52\]\[19\] _05265_ _05275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13514_ memory\[4\]\[29\] memory\[5\]\[29\] _05789_ _02903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14494_ _01533_ clknet_leaf_352_clk_i memory\[23\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_458 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11038__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13445_ memory\[54\]\[28\] memory\[55\]\[28\] _02312_ _02835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10835__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10657_ _05238_ _00365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_845 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13376_ _02167_ _02766_ _05756_ _02767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_3_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_261_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08305__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10588_ _05201_ _00333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12327_ memory\[46\]\[11\] memory\[47\]\[11\] _05907_ _06532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15115_ _00074_ clknet_leaf_34_clk_i memory\[42\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_110_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_192_Right_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15046_ _00005_ clknet_leaf_32_clk_i memory\[40\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09403__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12258_ _06325_ _06463_ _06464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_361_clk_i clknet_5_3__leaf_clk_i clknet_leaf_361_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_142_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12163__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11209_ _05531_ _00624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11210__I0 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12189_ memory\[30\]\[9\] memory\[31\]\[9\] _06193_ _06396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08040__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11465__I _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12070__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_376_clk_i clknet_5_12__leaf_clk_i clknet_leaf_376_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08975__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07717__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_108_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_92_57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08390__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08420_ _03762_ memory\[20\]\[5\] _04001_ _04007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13415__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08351_ _03970_ _01407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13510__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_110_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08142__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07302_ _03393_ _00935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08282_ _03760_ memory\[18\]\[4\] _03929_ _03934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09890__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_73_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07233_ _03349_ _00910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_314_clk_i clknet_5_11__leaf_clk_i clknet_leaf_314_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10745__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11729__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13121__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07164_ _03301_ _00889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07095_ _03263_ _00858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_329_clk_i clknet_5_10__leaf_clk_i clknet_leaf_329_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_160_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08014__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12154__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11201__I0 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07956__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11901__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13076__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09805_ memory\[3\]\[18\] _03180_ _04762_ _04771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_31_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input39_I we_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13329__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07997_ _03771_ _01252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06948_ _03166_ memory\[14\]\[13\] _03157_ _03167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09736_ _04612_ memory\[38\]\[18\] _04725_ _04734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13654__A1 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07708__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09667_ _04697_ _01996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06879_ _03110_ _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_97_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08618_ _04112_ _01532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09598_ _04610_ memory\[36\]\[17\] _04653_ _04661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08549_ _04075_ _01500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11968__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_46_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11560_ _05772_ _05774_ _05775_ _05776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_135_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10511_ _05035_ memory\[4\]\[14\] _05156_ _05161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11491_ memory\[6\]\[0\] memory\[7\]\[0\] _05706_ _05707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13230_ _02623_ _02624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10442_ _05124_ _00264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09633__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13161_ _02213_ _02555_ _02352_ _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA_clkbuf_2_0_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10373_ _05033_ memory\[47\]\[13\] _05084_ _05088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12112_ memory\[44\]\[8\] memory\[45\]\[8\] _06319_ _06320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13092_ memory\[46\]\[22\] memory\[47\]\[22\] _02487_ _02488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12145__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12043_ _05760_ _06251_ _06252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10390__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12696__A2 _02090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09561__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15802_ _00761_ clknet_leaf_26_clk_i net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08795__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13645__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_208_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13994_ _01033_ clknet_leaf_232_clk_i memory\[59\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15733_ _00692_ clknet_leaf_149_clk_i memory\[61\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12945_ _02341_ _02342_ _06866_ _02343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13206__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15664_ _00623_ clknet_leaf_144_clk_i memory\[5\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12876_ _06453_ _02274_ _02275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__11259__I0 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_103_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14615_ _01654_ clknet_leaf_79_clk_i memory\[26\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_103_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11827_ _05661_ _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_190_4036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08124__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15595_ _00554_ clknet_leaf_230_clk_i memory\[57\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11959__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14546_ _01585_ clknet_leaf_82_clk_i memory\[24\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11758_ _05741_ _05970_ _05971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_44_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08675__I1 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12620__A2 _06790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07003__I net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10709_ _05266_ _00389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14477_ _01516_ clknet_leaf_182_clk_i memory\[22\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11689_ _05741_ _05902_ _05903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_37_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13428_ _02371_ _02818_ _02373_ _02819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_148_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11431__I0 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13359_ memory\[24\]\[26\] memory\[25\]\[26\] memory\[26\]\[26\] memory\[27\]\[26\]
+ _02363_ _02502_ _02751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_80_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_23_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07874__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_149_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12136__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11396__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07920_ _03724_ _01222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15029_ _02068_ clknet_leaf_57_clk_i memory\[3\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08769__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07938__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07851_ _03160_ memory\[7\]\[11\] _03686_ _03688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_127_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07782_ _03651_ _01157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xinput2 address_i[1] net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_56_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09521_ _03183_ _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_91_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08363__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11742__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09452_ _04568_ _01910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10170__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08403_ _03997_ _01432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09383_ _04239_ memory\[33\]\[27\] _04524_ _04532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08334_ _03812_ memory\[18\]\[29\] _03951_ _03961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09863__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_253_clk_i clknet_5_24__leaf_clk_i clknet_leaf_253_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_188_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08265_ _03924_ _01367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07848__I _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_175_Left_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07216_ _03168_ _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_132_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08196_ _03810_ memory\[29\]\[28\] _03879_ _03888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09615__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07147_ _03194_ memory\[13\]\[22\] _03290_ _03293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_4_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_268_clk_i clknet_5_13__leaf_clk_i clknet_leaf_268_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_157_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_186_3949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07078_ _03197_ memory\[16\]\[23\] _03251_ _03255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12703__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07929__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_7_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_184_Left_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_22_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_87_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09504__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_206_clk_i clknet_5_31__leaf_clk_i clknet_leaf_206_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_173_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09719_ _04713_ _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10991_ _05037_ memory\[56\]\[15\] _05410_ _05416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08354__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13026__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_48_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12730_ memory\[36\]\[17\] memory\[37\]\[17\] _06447_ _02131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12661_ _06713_ _06856_ _06858_ _06860_ _06861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12865__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14400_ _01439_ clknet_leaf_352_clk_i memory\[20\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11612_ _05826_ _05827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_154_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12592_ memory\[38\]\[15\] memory\[39\]\[15\] _06728_ _06793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15380_ _00339_ clknet_leaf_155_clk_i memory\[50\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08657__I1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09854__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_193_Left_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14331_ _01370_ clknet_leaf_27_clk_i memory\[17\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_61_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11543_ _03117_ _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_9_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_53_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_61_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10385__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_491 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14262_ _01301_ clknet_leaf_138_clk_i memory\[15\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11474_ _05689_ _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_190_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12366__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13213_ _02319_ _02599_ _02606_ _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__13696__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11413__I0 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10425_ _05115_ _00256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14193_ _01232_ clknet_leaf_117_clk_i memory\[19\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09082__I1 memory\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09973__I _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07694__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13144_ _02538_ _02539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10356_ _05016_ memory\[47\]\[5\] _05073_ _05079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13075_ memory\[14\]\[22\] memory\[15\]\[22\] _02193_ _02471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10912__I _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10287_ _05033_ memory\[46\]\[13\] _05027_ _05034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12026_ _06028_ _06234_ _05722_ _06235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_100_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_359_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13977_ _01016_ clknet_leaf_382_clk_i memory\[49\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15716_ _00675_ clknet_leaf_310_clk_i memory\[61\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12928_ _06851_ _02325_ _02326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10152__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15647_ _00606_ clknet_leaf_367_clk_i memory\[5\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12775__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12859_ _06848_ _02257_ _06707_ _02258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__13477__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_173_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_411_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08648__I1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15578_ _00537_ clknet_leaf_373_clk_i memory\[56\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14529_ _01568_ clknet_leaf_354_clk_i memory\[24\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07320__I1 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08050_ _03807_ _01269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_153_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07001_ _03206_ memory\[14\]\[26\] _03188_ _03207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12357__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11404__I0 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_168_3613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09073__I1 memory\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07084__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12109__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10822__I _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08952_ _04216_ memory\[27\]\[16\] _04297_ _04304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07109__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07903_ _03715_ _01214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08883_ _04267_ _01642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_181_3857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07834_ _03135_ memory\[7\]\[3\] _03675_ _03679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06948__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07765_ _03642_ _01149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09504_ _04602_ memory\[35\]\[13\] _04596_ _04603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07696_ _03132_ memory\[63\]\[2\] _03603_ _03606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10143__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09435_ _04559_ _01902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_83_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_192_clk_i clknet_5_29__leaf_clk_i clknet_leaf_192_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_149_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09366_ _04222_ memory\[33\]\[19\] _04513_ _04523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_81_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08317_ _03952_ _01391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09297_ _04486_ _01837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_394 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__I1 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08248_ _03793_ memory\[17\]\[20\] _03915_ _03916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12348__A1 _06507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08179_ _03856_ _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_15_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10210_ _04986_ _00170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11190_ _05521_ _00615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_130_clk_i clknet_5_22__leaf_clk_i clknet_leaf_130_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_101_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10141_ _04606_ memory\[44\]\[15\] _04944_ _04950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_89_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10072_ _04913_ _00105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08575__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13900_ _00939_ clknet_leaf_214_clk_i memory\[11\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_145_clk_i clknet_5_22__leaf_clk_i clknet_leaf_145_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14880_ _01919_ clknet_leaf_420_clk_i memory\[35\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_360_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_921 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13831_ _00870_ clknet_leaf_202_clk_i memory\[13\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_67_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11563__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10974_ _05020_ memory\[56\]\[7\] _05399_ _05407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13762_ _00801_ clknet_leaf_281_clk_i memory\[14\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_63_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15501_ _00460_ clknet_leaf_240_clk_i memory\[54\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_63_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12713_ _06831_ _02109_ _02111_ _02113_ _02114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_100_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13693_ _03077_ _00764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_100_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07550__I1 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15432_ _00391_ clknet_leaf_296_clk_i memory\[52\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12644_ _05652_ _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_80_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13623__I1 net63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12587__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12608__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15363_ _00322_ clknet_leaf_335_clk_i memory\[50\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12575_ _06775_ _06776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_182_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11004__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14314_ _01353_ clknet_leaf_207_clk_i memory\[17\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11526_ _05669_ _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15294_ _00253_ clknet_leaf_347_clk_i memory\[48\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12339__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11457_ _05668_ _05672_ _05673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14245_ _01284_ clknet_leaf_276_clk_i memory\[15\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09409__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10408_ _05068_ memory\[47\]\[30\] _05072_ _05106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14176_ _01215_ clknet_leaf_342_clk_i memory\[19\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_78_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08313__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11388_ _05626_ _00708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13439__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12343__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13127_ _02163_ _02517_ _02519_ _02521_ _02522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10339_ _05068_ memory\[46\]\[30\] _05005_ _05069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_163_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_163_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12198__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13058_ memory\[52\]\[22\] memory\[53\]\[22\] _06832_ _02454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12009_ _06217_ _06218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10373__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09144__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08318__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11473__I _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_105_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07550_ memory\[59\]\[31\] _03373_ _03492_ _03527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08983__S _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07481_ _03489_ _01018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09220_ _04212_ memory\[31\]\[14\] _04441_ _04446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07599__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08782__I _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09151_ _04409_ _01768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_90_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_20_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08102_ _03837_ _01291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09082_ _04210_ memory\[2\]\[13\] _04369_ _04373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08033_ _03190_ _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_135_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_135_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07057__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09319__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12750__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09984_ _04585_ memory\[42\]\[5\] _04861_ _04867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_clk_i clknet_5_16__leaf_clk_i clknet_leaf_62_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08935_ _04199_ memory\[27\]\[8\] _04286_ _04295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08866_ _04258_ _01634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10364__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input21_I data_i[22] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07817_ _03669_ _01174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08797_ _03171_ _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08309__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_84_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_77_clk_i clknet_5_17__leaf_clk_i clknet_leaf_77_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07748_ _03209_ memory\[63\]\[27\] _03625_ _03633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_28_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08893__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10116__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10667__I1 _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07679_ _03596_ _01109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07532__I1 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09788__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09418_ _04206_ memory\[34\]\[11\] _04549_ _04551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10690_ _05256_ _00380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12569__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09349_ _04514_ _01861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_307_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12360_ _06563_ _06564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_105_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11311_ memory\[61\]\[5\] _03140_ _05580_ _05586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_15_clk_i clknet_5_5__leaf_clk_i clknet_leaf_15_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12291_ _06276_ _06495_ _06001_ _06496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10663__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14030_ _01069_ clknet_leaf_170_clk_i memory\[0\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07048__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11242_ _03319_ memory\[60\]\[5\] _05543_ _05549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12592__I1 memory\[39\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11173_ _05512_ _00607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_56_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09028__I _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_56_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07972__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10124_ _04589_ memory\[44\]\[7\] _04933_ _04941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08548__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10055_ _04904_ _00097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14932_ _01971_ clknet_leaf_12_clk_i memory\[36\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07220__I0 memory\[39\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11507__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14863_ _01902_ clknet_leaf_63_clk_i memory\[34\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13814_ _00853_ clknet_leaf_110_clk_i memory\[16\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14794_ _01833_ clknet_leaf_44_clk_i memory\[32\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13745_ _03104_ _00789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10658__I1 _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10957_ _05397_ _00506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08476__A2 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08720__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07523__I1 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09698__I _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13214__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11480__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_139_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13676_ _02494_ _03058_ _03060_ _03062_ _03063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_10888_ _05360_ _00474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15415_ _00374_ clknet_leaf_382_clk_i memory\[51\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12627_ _03120_ _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_156_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_5_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15346_ _00305_ clknet_leaf_145_clk_i memory\[4\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12558_ _06759_ _00745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07011__I net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12980__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11783__A2 _05965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11509_ _05691_ _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10573__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15277_ _00236_ clknet_leaf_277_clk_i memory\[47\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12489_ _06276_ _06689_ _06690_ _06691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_151_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09139__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14228_ _01267_ clknet_leaf_114_clk_i memory\[12\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08043__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13169__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11468__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14159_ _01198_ clknet_leaf_218_clk_i memory\[7\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_130_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10594__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07882__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_130_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06981_ _03191_ memory\[14\]\[21\] _03188_ _03192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08720_ _03789_ memory\[24\]\[18\] _04157_ _04166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10346__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08651_ _04129_ _01548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07211__I0 memory\[39\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07602_ _03555_ _01073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_256_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08582_ _04092_ _01516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12799__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09602__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07533_ _03518_ _01041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_176_3767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_146_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07464_ memory\[49\]\[23\] _03357_ _03477_ _03481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08218__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07122__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09203_ _04195_ memory\[31\]\[6\] _04430_ _04437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07395_ _03442_ _00979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12963__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09134_ _04400_ _01760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08017__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09065_ _04193_ memory\[2\]\[5\] _04358_ _04364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_4_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08016_ _03784_ _01258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09049__S _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_38_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08888__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10585__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09967_ _04857_ _00056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08918_ _04285_ _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12203__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09898_ _04635_ memory\[40\]\[29\] _04811_ _04821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_51_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_14__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08849_ net72 _03855_ _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08950__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11860_ memory\[60\]\[5\] memory\[61\]\[5\] _05656_ _06071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13542__B _02928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10811_ _05062_ memory\[53\]\[27\] _05312_ _05320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11791_ memory\[56\]\[4\] memory\[57\]\[4\] memory\[58\]\[4\] memory\[59\]\[4\] _05670_
+ _05671_ _06003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10658__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13034__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13530_ _02918_ _02919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06935__I _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10742_ _05283_ _00405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08128__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07032__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13461_ _05772_ _02850_ _05775_ _02851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_138_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10673_ memory\[51\]\[26\] _03205_ _05240_ _05247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12873__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_173_Right_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15200_ _00159_ clknet_leaf_423_clk_i memory\[45\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12412_ _06615_ _06616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_129_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_11_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_97_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13392_ memory\[0\]\[27\] memory\[1\]\[27\] memory\[2\]\[27\] memory\[3\]\[27\] _05784_
+ _03226_ _02783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15131_ _00090_ clknet_leaf_441_clk_i memory\[42\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12343_ _06480_ _06547_ _06482_ _06548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_58_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_58_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12274_ _05752_ _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15062_ _00021_ clknet_leaf_7_clk_i memory\[40\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12714__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13062__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14013_ _01052_ clknet_leaf_371_clk_i memory\[0\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11225_ _05539_ _00632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08798__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11156_ _03369_ memory\[58\]\[29\] _05493_ _05503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10107_ _04931_ _00122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11087_ _05466_ _00567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_175_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14915_ _01954_ clknet_leaf_432_clk_i memory\[36\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10038_ _04639_ memory\[42\]\[31\] _04860_ _04895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_37_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14846_ _01885_ clknet_leaf_424_clk_i memory\[34\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09422__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_19_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10568__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14777_ _01816_ clknet_leaf_60_clk_i memory\[31\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11989_ _05914_ _06192_ _06196_ _06198_ _06199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_105_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_193_4078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13728_ _03095_ _00781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10500__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_154_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13659_ memory\[32\]\[31\] memory\[33\]\[31\] memory\[34\]\[31\] memory\[35\]\[31\]
+ _05670_ _05671_ _03046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12628__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_140_Right_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_26_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07180_ memory\[39\]\[2\] _03313_ _03309_ _03314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_171_3675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15329_ _00288_ clknet_leaf_340_clk_i memory\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07680__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12705__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09821_ _04779_ _02068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08501__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13119__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12023__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09752_ _04742_ _02036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06964_ _03178_ memory\[14\]\[17\] _03157_ _03179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09185__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08703_ _04145_ _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_6_Left_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06895_ _03111_ memory\[14\]\[0\] _03126_ _03127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09683_ _04627_ memory\[37\]\[25\] _04700_ _04706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11862__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08634_ _04120_ _01540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06956__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_94_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_167_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08565_ _04083_ _01508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10478__S _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13433__A2 _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12867__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07516_ _03509_ _01033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08496_ _03770_ memory\[21\]\[9\] _04037_ _04047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10277__I _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07447_ memory\[49\]\[15\] _03340_ _03466_ _03472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07787__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13197__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07378_ _03433_ _00971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08999__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11610__B _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09117_ _04245_ memory\[2\]\[30\] _04357_ _04391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08612__A2 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11102__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09048_ _04354_ _01720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13744__I0 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10558__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11010_ _05056_ memory\[56\]\[24\] _05421_ _05426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_53_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09507__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output52_I net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12961_ memory\[28\]\[20\] memory\[29\]\[20\] _06604_ _02359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14700_ _01739_ clknet_leaf_172_clk_i memory\[2\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08923__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11912_ _05914_ _06118_ _06120_ _06122_ _06123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15680_ _00639_ clknet_leaf_323_clk_i memory\[60\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11683__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12892_ _06603_ _02286_ _02288_ _02290_ _02291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_158_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_99_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12307__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13272__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14631_ _01670_ clknet_leaf_179_clk_i memory\[27\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11843_ memory\[30\]\[4\] memory\[31\]\[4\] _05773_ _06055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10388__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_16_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14562_ _01601_ clknet_leaf_408_clk_i memory\[25\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11774_ _05914_ _05982_ _05984_ _05986_ _05987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_99_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13513_ _02302_ _02894_ _02901_ _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_10725_ _05274_ _00397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14493_ _01532_ clknet_leaf_358_clk_i memory\[23\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13444_ _02833_ _02834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10656_ memory\[51\]\[18\] _03180_ _05229_ _05238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12935__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_204_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13375_ memory\[62\]\[27\] memory\[63\]\[27\] _02448_ _02766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10587_ _05043_ memory\[50\]\[18\] _05192_ _05201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10797__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15114_ _00073_ clknet_leaf_21_clk_i memory\[42\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12326_ _06530_ _06531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_121_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_110_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11947__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15045_ _00004_ clknet_leaf_431_clk_i memory\[40\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12257_ memory\[40\]\[10\] memory\[41\]\[10\] memory\[42\]\[10\] memory\[43\]\[10\]
+ _06186_ _06326_ _06463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_82_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13360__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11208_ _03353_ memory\[5\]\[21\] _05529_ _05531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12188_ _06394_ _06395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_43_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_79_Left_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11139_ _05494_ _00591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09167__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11674__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09152__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_125_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07342__A2 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14829_ _01868_ clknet_leaf_51_clk_i memory\[33\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13415__A2 _02805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08350_ _03760_ memory\[1\]\[4\] _03965_ _03970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_173_3704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08991__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07301_ memory\[11\]\[12\] _03334_ _03390_ _03393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_88_Left_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08281_ _03933_ _01374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13179__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07232_ memory\[39\]\[19\] _03348_ _03330_ _03349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07400__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12926__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07163_ _03218_ memory\[13\]\[30\] _03267_ _03301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12018__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10788__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07653__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07094_ _03221_ memory\[16\]\[31\] _03228_ _03263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10761__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09327__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_97_Left_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08231__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_406_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09804_ _04770_ _02060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_31_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10960__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07996_ _03770_ memory\[12\]\[9\] _03752_ _03771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09158__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08030__I _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09735_ _04733_ _02028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06947_ _03165_ _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08905__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11665__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09666_ _04610_ memory\[37\]\[17\] _04689_ _04697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06878_ net7 _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_59_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10712__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08617_ memory\[23\]\[1\] _03311_ _04110_ _04112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_153_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09597_ _04660_ _01963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09997__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10001__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08548_ _03754_ memory\[22\]\[1\] _04073_ _04075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07097__A1 _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12090__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08479_ _04038_ _01467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_46_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_421_clk_i clknet_5_0__leaf_clk_i clknet_leaf_421_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13312__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10510_ _05160_ _00296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07892__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11490_ _05661_ _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08406__S _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10441_ _05033_ memory\[48\]\[13\] _05120_ _05124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13590__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08205__I _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13160_ memory\[46\]\[23\] memory\[47\]\[23\] _02487_ _02555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10372_ _05087_ _00231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_436_clk_i clknet_5_0__leaf_clk_i clknet_leaf_436_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_60_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13717__I0 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12111_ _05677_ _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13091_ _05701_ _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10671__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_78_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09237__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09397__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12042_ memory\[40\]\[7\] memory\[41\]\[7\] memory\[42\]\[7\] memory\[43\]\[7\] _06186_
+ _05762_ _06251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_1_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_40_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15801_ _00760_ clknet_leaf_62_clk_i net61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13993_ _01032_ clknet_leaf_233_clk_i memory\[59\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15732_ _00691_ clknet_leaf_162_clk_i memory\[61\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11656__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12944_ memory\[38\]\[20\] memory\[39\]\[20\] _06728_ _02342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10703__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15663_ _00622_ clknet_leaf_250_clk_i memory\[5\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12875_ memory\[32\]\[19\] memory\[33\]\[19\] memory\[34\]\[19\] memory\[35\]\[19\]
+ _02205_ _06454_ _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
Xclkbuf_5_8__f_clk_i clknet_2_1_0_clk_i clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_185_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14614_ _01653_ clknet_leaf_82_clk_i memory\[26\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_103_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11826_ _06037_ _06038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_190_4026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_103_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15594_ _00553_ clknet_leaf_231_clk_i memory\[57\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_190_4037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09321__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14545_ _01584_ clknet_leaf_93_clk_i memory\[24\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11757_ memory\[32\]\[3\] memory\[33\]\[3\] memory\[34\]\[3\] memory\[35\]\[3\] _05742_
+ _05743_ _05970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10846__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12620__A3 _06805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10708_ _05026_ memory\[52\]\[10\] _05265_ _05266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08316__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14476_ _01515_ clknet_leaf_174_clk_i memory\[22\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11688_ memory\[32\]\[2\] memory\[33\]\[2\] memory\[34\]\[2\] memory\[35\]\[2\] _05742_
+ _05743_ _05902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_183_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12908__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_355_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13427_ memory\[22\]\[27\] memory\[23\]\[27\] _05754_ _02818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10639_ _05217_ _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_113_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_148_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_84_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13358_ _02498_ _02749_ _05665_ _02750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11677__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13708__I0 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12309_ _06155_ _06509_ _06511_ _06513_ _06514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__10581__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13289_ _02216_ _02681_ _02682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_149_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15028_ _02067_ clknet_leaf_57_clk_i memory\[3\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_18_Right_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11195__I0 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11476__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07850_ _03687_ _01189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_127_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07890__S _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_127_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07781_ _03156_ memory\[6\]\[10\] _03650_ _03651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput3 address_i[2] net3 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_78_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09520_ _04613_ _01933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08785__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11647__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11742__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09451_ _04239_ memory\[34\]\[27\] _04560_ _04568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08402_ _03812_ memory\[1\]\[29\] _03987_ _03997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09382_ _04531_ _01877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_27_Right_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08333_ _03960_ _01399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_145_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08264_ _03810_ memory\[17\]\[28\] _03915_ _03924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07874__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07130__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12256__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07215_ _03337_ _00904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12971__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08195_ _03887_ _01334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_41_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07146_ _03292_ _00880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13572__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07626__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11587__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07077_ _03254_ _00849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12770__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_36_Right_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13324__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09057__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11886__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07979_ _03759_ _01246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09718_ _04724_ _02020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10990_ _05415_ _00521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07305__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09649_ _04593_ memory\[37\]\[9\] _04678_ _04688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_48_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Right_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13106__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12660_ _06720_ _06859_ _06860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_65_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_360_clk_i clknet_5_3__leaf_clk_i clknet_leaf_360_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09303__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11611_ memory\[12\]\[1\] memory\[13\]\[1\] _05716_ _05826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11110__I0 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12591_ _06791_ _06792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_110_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14330_ _01369_ clknet_leaf_26_clk_i memory\[17\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07865__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06943__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11542_ _05753_ _05755_ _05757_ _05758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_37_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11810__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_61_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07040__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14261_ _01300_ clknet_leaf_112_clk_i memory\[15\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11473_ _03117_ _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xclkbuf_leaf_375_clk_i clknet_5_9__leaf_clk_i clknet_leaf_375_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13212_ _05768_ _02601_ _02603_ _02605_ _02606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07975__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10424_ _05016_ memory\[48\]\[5\] _05109_ _05115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07617__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14192_ _01231_ clknet_leaf_103_clk_i memory\[19\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_54_Right_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_21_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13143_ memory\[12\]\[23\] memory\[13\]\[23\] _06714_ _02538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08290__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10355_ _05078_ _00223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13315__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12749__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13074_ _02469_ _02470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10286_ _03165_ _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_40_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12025_ memory\[14\]\[7\] memory\[15\]\[7\] _05720_ _06234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_144_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_144_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_313_clk_i clknet_5_11__leaf_clk_i clknet_leaf_313_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_161_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11629__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_105_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_189_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_161_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_105_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13976_ _01015_ clknet_leaf_382_clk_i memory\[49\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_63_Right_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15715_ _00674_ clknet_leaf_322_clk_i memory\[61\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12927_ memory\[0\]\[20\] memory\[1\]\[20\] memory\[2\]\[20\] memory\[3\]\[20\] _06709_
+ _06779_ _02325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_122_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15646_ _00605_ clknet_leaf_369_clk_i memory\[5\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12858_ memory\[6\]\[19\] memory\[7\]\[19\] _06431_ _02257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_328_clk_i clknet_5_10__leaf_clk_i clknet_leaf_328_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_158_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13477__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09430__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11809_ memory\[0\]\[4\] memory\[1\]\[4\] memory\[2\]\[4\] memory\[3\]\[4\] _06020_
+ _03748_ _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_15577_ _00536_ clknet_leaf_271_clk_i memory\[56\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12789_ _06851_ _02188_ _02189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_173_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11801__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14528_ _01567_ clknet_leaf_354_clk_i memory\[24\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08046__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12791__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14459_ _01498_ clknet_leaf_0_clk_i memory\[21\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07000_ _03205_ _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XPHY_EDGE_ROW_72_Right_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13554__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_101_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12804__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13306__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08951_ _04303_ _01674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11168__I0 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07902_ _03135_ memory\[19\]\[3\] _03711_ _03715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08882_ _04214_ memory\[26\]\[15\] _04261_ _04267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_181_3858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09605__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13635__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07833_ _03678_ _01181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_81_Right_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12031__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07764_ _03132_ memory\[6\]\[2\] _03639_ _03642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09503_ _03165_ _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_56_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12293__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07695_ _03605_ _01116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_26_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09434_ _04222_ memory\[34\]\[19\] _04549_ _04559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06964__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_136_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12045__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11479__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10486__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09365_ _04522_ _01869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_23_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_43_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08316_ _03793_ memory\[18\]\[20\] _03951_ _03952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_23_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09296_ _04220_ memory\[32\]\[18\] _04477_ _04486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Right_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_16_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08247_ _03892_ _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_166_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07795__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12348__A2 _06522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12979__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08178_ _03878_ _01326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_166_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07129_ _03283_ _00872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12206__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11110__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10140_ _04949_ _00137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_89_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08024__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10071_ _04604_ memory\[43\]\[14\] _04908_ _04913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_89_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_303_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13830_ _00869_ clknet_leaf_201_clk_i memory\[13\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06938__I net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_26__f_clk_i clknet_2_3_0_clk_i clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13761_ _00800_ clknet_leaf_280_clk_i memory\[14\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12284__A1 _06427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10973_ _05406_ _00513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15500_ _00459_ clknet_leaf_290_clk_i memory\[54\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12712_ _06838_ _02112_ _02113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_63_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13692_ _03311_ memory\[9\]\[1\] _03075_ _03077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_100_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15431_ _00390_ clknet_leaf_295_clk_i memory\[52\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13280__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12036__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12675__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10396__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12643_ _06411_ _06830_ _06842_ _06843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_80_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_80_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12587__A2 _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15362_ _00321_ clknet_leaf_314_clk_i memory\[50\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07838__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12574_ memory\[4\]\[15\] memory\[5\]\[15\] _06156_ _06775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14313_ _01352_ clknet_leaf_208_clk_i memory\[17\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11525_ _05667_ _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_15293_ _00252_ clknet_leaf_345_clk_i memory\[48\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_29_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_68_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14244_ _01283_ clknet_leaf_276_clk_i memory\[15\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11456_ memory\[56\]\[0\] memory\[57\]\[0\] memory\[58\]\[0\] memory\[59\]\[0\] _05670_
+ _05671_ _05672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_80_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11398__I0 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_3__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10407_ _05105_ _00248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14175_ _01214_ clknet_leaf_357_clk_i memory\[19\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11387_ _03327_ memory\[62\]\[9\] _05616_ _05626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_78_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11020__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13126_ _02170_ _02520_ _02521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10338_ _03217_ _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_178_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08015__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12198__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13057_ _02163_ _02447_ _02450_ _02452_ _02453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10269_ _05021_ _00194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_252_clk_i clknet_5_25__leaf_clk_i clknet_leaf_252_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12008_ memory\[52\]\[7\] memory\[53\]\[7\] _06143_ _06217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09763__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13147__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_187_Right_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12786__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13959_ _00998_ clknet_leaf_295_clk_i memory\[49\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_267_clk_i clknet_5_13__leaf_clk_i clknet_leaf_267_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_124_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07480_ memory\[49\]\[31\] _03373_ _03454_ _03489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09160__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15629_ _00588_ clknet_leaf_228_clk_i memory\[58\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09818__I1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09150_ _04210_ memory\[30\]\[13\] _04405_ _04409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08101_ _03785_ memory\[15\]\[16\] _03830_ _03837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09081_ _04372_ _01735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_12_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_15_Left_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13527__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13410__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08032_ _03795_ _01263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_135_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_135_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_252_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_205_clk_i clknet_5_31__leaf_clk_i clknet_leaf_205_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_3_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_163_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08254__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09983_ _04866_ _00063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_1339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08006__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08934_ _04294_ _01666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09335__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13365__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08865_ _04197_ memory\[26\]\[7\] _04250_ _04258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_24_Left_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_93_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07816_ _03209_ memory\[6\]\[27\] _03661_ _03669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08796_ _04213_ _01609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input14_I data_i[16] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07747_ _03632_ _01141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_154_Right_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07678_ _03206_ memory\[10\]\[26\] _03589_ _03596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_0_Right_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09417_ _04550_ _01893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_164_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09348_ _04203_ memory\[33\]\[10\] _04513_ _04514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_33_Left_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10944__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09279_ _04465_ _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_7_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11310_ _05585_ _00671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12290_ memory\[62\]\[11\] memory\[63\]\[11\] _05868_ _06495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08414__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08245__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11241_ _05548_ _00639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10052__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11172_ _03317_ memory\[5\]\[4\] _05507_ _05512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_56_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11775__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10123_ _04940_ _00129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13377__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_42_Left_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09245__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09745__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10054_ _04587_ memory\[43\]\[6\] _04897_ _04904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14931_ _01970_ clknet_leaf_73_clk_i memory\[36\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07220__I1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14862_ _01901_ clknet_leaf_63_clk_i memory\[34\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13813_ _00852_ clknet_leaf_114_clk_i memory\[16\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14793_ _01832_ clknet_leaf_43_clk_i memory\[32\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_121_Right_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_98_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13744_ _03363_ memory\[9\]\[26\] _03097_ _03104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10956_ memory\[55\]\[31\] _03220_ _05362_ _05397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13675_ _02501_ _03061_ _03062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_183_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10887_ _05070_ memory\[54\]\[31\] _05325_ _05360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_139_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_51_Left_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_38_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15414_ _00373_ clknet_leaf_42_clk_i memory\[51\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12626_ _06276_ _06825_ _06690_ _06826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_183_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15345_ _00304_ clknet_leaf_144_clk_i memory\[4\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08484__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10854__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12557_ _06758_ net45 _06491_ _06759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_117_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13509__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11508_ _05689_ _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08324__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11783__A3 _05980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15276_ _00235_ clknet_leaf_271_clk_i memory\[47\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12488_ _05664_ _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_53_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_0_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09189__A1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14227_ _01266_ clknet_leaf_118_clk_i memory\[12\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11439_ _03120_ _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11615__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09984__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14158_ _01197_ clknet_leaf_219_clk_i memory\[7\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_130_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_60_Left_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_191_clk_i clknet_5_29__leaf_clk_i clknet_leaf_191_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13109_ _02494_ _02497_ _02500_ _02504_ _02505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_130_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06980_ _03190_ _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_14089_ _01128_ clknet_leaf_223_clk_i memory\[63\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07962__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input6_I address_i[5] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09736__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12496__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11484__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08650_ memory\[23\]\[17\] _03344_ _04121_ _04129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07211__I1 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_179_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07601_ _03194_ memory\[0\]\[22\] _03552_ _03555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08581_ _03787_ memory\[22\]\[17\] _04084_ _04092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13405__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07532_ memory\[59\]\[22\] _03355_ _03515_ _03518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13540__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07463_ _03480_ _01009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09202_ _04436_ _01792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_63_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07394_ _03200_ memory\[8\]\[24\] _03437_ _03442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09133_ _04193_ memory\[30\]\[5\] _04394_ _04400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07278__I1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_144_clk_i clknet_5_22__leaf_clk_i clknet_leaf_144_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09064_ _04363_ _01727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08015_ _03783_ memory\[12\]\[15\] _03773_ _03784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08227__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10034__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08033__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_38_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_159_clk_i clknet_5_24__leaf_clk_i clknet_leaf_159_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13359__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09966_ _04635_ memory\[41\]\[29\] _04847_ _04857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09065__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08917_ _03376_ _03855_ _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_09897_ _04820_ _00023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_51_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08848_ _04248_ _01626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08779_ _04201_ memory\[25\]\[9\] _04183_ _04202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10810_ _05319_ _00437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_170_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11790_ _05660_ _06000_ _06001_ _06002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_68_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07313__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10741_ _05060_ memory\[52\]\[26\] _05276_ _05283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13460_ memory\[14\]\[28\] memory\[15\]\[28\] _05773_ _02850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12098__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10672_ _05246_ _00372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12411_ memory\[20\]\[12\] memory\[21\]\[12\] _06477_ _06615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08466__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07269__I1 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13391_ _05752_ _02781_ _05791_ _02782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_11_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11845__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_97_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13050__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_97_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15130_ _00089_ clknet_leaf_441_clk_i memory\[42\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12342_ memory\[22\]\[11\] memory\[23\]\[11\] _06062_ _06547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06951__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08144__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11569__I _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_58_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08218__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15061_ _00020_ clknet_leaf_9_clk_i memory\[40\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12273_ _06478_ _06479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_82_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_148_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14012_ _01051_ clknet_leaf_371_clk_i memory\[0\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09966__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11224_ _03369_ memory\[5\]\[29\] _05529_ _05539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12714__A2 _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11155_ _05502_ _00599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07441__I1 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10106_ _04639_ memory\[43\]\[31\] _04896_ _04931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11086_ _05064_ memory\[57\]\[28\] _05457_ _05466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14914_ _01953_ clknet_leaf_432_clk_i memory\[36\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10037_ _04894_ _00089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_200_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09703__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14845_ _01884_ clknet_leaf_429_clk_i memory\[34\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06952__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14776_ _01815_ clknet_leaf_60_clk_i memory\[31\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_158_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11988_ _05921_ _06197_ _06198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13727_ _03346_ memory\[9\]\[18\] _03086_ _03095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_193_4079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12650__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10939_ _05388_ _00497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_184_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13658_ _05660_ _03044_ _05708_ _03045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12089__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_61_clk_i clknet_5_17__leaf_clk_i clknet_leaf_61_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_27_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12609_ memory\[24\]\[15\] memory\[25\]\[15\] memory\[26\]\[15\] memory\[27\]\[15\]
+ _06472_ _06611_ _06810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_170_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13589_ _05777_ _02976_ _02977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15328_ _00287_ clknet_leaf_340_clk_i memory\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_30_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15259_ _00218_ clknet_leaf_392_clk_i memory\[46\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08989__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_76_clk_i clknet_5_16__leaf_clk_i clknet_leaf_76_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10016__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09820_ memory\[3\]\[25\] _03202_ _04773_ _04779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08788__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07432__I1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09709__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09751_ _04627_ memory\[38\]\[25\] _04736_ _04742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06963_ _03177_ _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_33_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_33_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08702_ _04156_ _01572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09682_ _04705_ _02003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_06894_ _03125_ _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09613__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08633_ memory\[23\]\[9\] _03327_ _04110_ _04120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_178_3808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13643__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10759__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_14_clk_i clknet_5_5__leaf_clk_i clknet_leaf_14_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08564_ _03770_ memory\[22\]\[9\] _04073_ _04083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08229__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13433__A3 _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07515_ memory\[59\]\[14\] _03338_ _03504_ _03509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12974__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08495_ _04046_ _01475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12641__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_146_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_clk_i clknet_5_4__leaf_clk_i clknet_leaf_29_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07446_ _03471_ _01001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_402_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10494__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07377_ _03175_ memory\[8\]\[16\] _03426_ _03433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09116_ _04390_ _01752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_107_Left_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_103_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11389__I _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09047_ _04243_ memory\[28\]\[29\] _04344_ _04354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_142_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08899__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10007__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09948__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_70_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09949_ _04848_ _00047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09325__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12960_ _03224_ _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XPHY_EDGE_ROW_116_Left_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output45_I net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11911_ _05921_ _06121_ _06122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_12891_ _06610_ _02289_ _02290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10669__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14630_ _01669_ clknet_leaf_179_clk_i memory\[27\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12307__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11842_ _06053_ _06054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__06946__I net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14561_ _01600_ clknet_leaf_414_clk_i memory\[25\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11773_ _05921_ _05985_ _05986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08687__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_74_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12483__I1 net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10494__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07978__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13512_ _05715_ _02896_ _02898_ _02900_ _02901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10724_ _05043_ memory\[52\]\[18\] _05265_ _05274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14492_ _01531_ clknet_leaf_362_clk_i memory\[23\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08439__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13443_ memory\[52\]\[28\] memory\[53\]\[28\] _05716_ _02833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10655_ _05237_ _00364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_180_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13374_ _02764_ _02765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_152_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07111__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10586_ _05200_ _00332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15113_ _00072_ clknet_leaf_25_clk_i memory\[42\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12325_ memory\[44\]\[11\] memory\[45\]\[11\] _06319_ _06530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_299_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15044_ _00003_ clknet_leaf_442_clk_i memory\[40\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09939__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_110_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12256_ _06322_ _06460_ _06461_ _06462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08602__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11207_ _05530_ _00623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12187_ memory\[28\]\[9\] memory\[29\]\[9\] _05915_ _06394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11138_ _03350_ memory\[58\]\[20\] _05493_ _05494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11069_ _05434_ _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_351_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10579__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14828_ _01867_ clknet_leaf_52_clk_i memory\[33\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08049__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09232__I _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12794__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14759_ _01798_ clknet_leaf_132_clk_i memory\[31\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07300_ _03392_ _00934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07888__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_59_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_665 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08280_ _03758_ memory\[18\]\[3\] _03929_ _03933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07350__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13689__I _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07231_ _03183_ _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11809__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11203__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12926__A2 _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07162_ _03300_ _00888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07093_ _03262_ _00857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08602__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07128__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09803_ memory\[3\]\[17\] _03177_ _04762_ _04770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07995_ _03152_ _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09734_ _04610_ memory\[38\]\[17\] _04725_ _04733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06946_ net11 _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__09343__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09665_ _04696_ _01995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12862__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08616_ _04111_ _01531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_136_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09596_ _04608_ memory\[36\]\[16\] _04653_ _04660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08547_ _04074_ _01499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10476__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07097__A2 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08478_ _03746_ memory\[21\]\[0\] _04037_ _04038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_46_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07429_ _03462_ _00993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_674 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_169_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_163_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10440_ _05123_ _00263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09094__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08841__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10952__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10371_ _05031_ memory\[47\]\[12\] _05084_ _05087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12110_ _05675_ _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08422__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_62_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13090_ _02485_ _02486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12041_ _05753_ _06249_ _05757_ _06250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_40_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07038__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10400__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15800_ _00759_ clknet_leaf_59_clk_i net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13992_ _01031_ clknet_leaf_233_clk_i memory\[59\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09253__S _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15731_ _00690_ clknet_leaf_148_clk_i memory\[61\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12943_ _05659_ _02341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12853__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06907__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15662_ _00621_ clknet_leaf_252_clk_i memory\[5\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12874_ _06450_ _02272_ _06866_ _02273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_87_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07580__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14613_ _01652_ clknet_leaf_81_clk_i memory\[26\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11825_ memory\[36\]\[4\] memory\[37\]\[4\] _05733_ _06037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10198__I _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15593_ _00552_ clknet_leaf_233_clk_i memory\[57\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_103_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_103_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14544_ _01583_ clknet_leaf_92_clk_i memory\[24\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11756_ _05736_ _05968_ _05739_ _05969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_83_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_120_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12620__A4 _06820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10707_ _05253_ _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14475_ _01514_ clknet_leaf_197_clk_i memory\[22\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11687_ _05736_ _05900_ _05739_ _05901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13426_ _02816_ _02817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_148_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10638_ _05228_ _00356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13030__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11958__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13357_ memory\[30\]\[26\] memory\[31\]\[26\] _05737_ _02749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10862__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08832__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10569_ _05191_ _00324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_11_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11592__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12308_ _06162_ _06512_ _06513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09428__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08332__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13288_ memory\[40\]\[25\] memory\[41\]\[25\] memory\[42\]\[25\] memory\[43\]\[25\]
+ _06875_ _02217_ _02681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__12362__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15027_ _02066_ clknet_leaf_139_clk_i memory\[3\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12239_ _03304_ _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_166_3564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10942__I1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07780_ _03638_ _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13097__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput4 address_i[3] net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_155_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08899__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11706__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12844__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11492__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09450_ _04567_ _01909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10102__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07571__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08401_ _03996_ _01431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09381_ _04237_ memory\[33\]\[26\] _04524_ _04531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08332_ _03810_ memory\[18\]\[28\] _03951_ _03960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10458__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_15_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08507__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08263_ _03923_ _01366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_62_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07214_ memory\[39\]\[13\] _03336_ _03330_ _03337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09076__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08194_ _03808_ memory\[29\]\[27\] _03879_ _03887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07210__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07145_ _03191_ memory\[13\]\[21\] _03290_ _03292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08823__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11583__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07076_ _03194_ memory\[16\]\[22\] _03251_ _03254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_22_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_7_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_7_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07978_ _03758_ memory\[12\]\[3\] _03752_ _03759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09073__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09717_ _04593_ memory\[38\]\[9\] _04714_ _04724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06929_ net38 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_87_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_87_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11108__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_247_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10697__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09648_ _04687_ _01987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_48_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09801__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09579_ _04591_ memory\[36\]\[8\] _04642_ _04651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11610_ _05700_ _05820_ _05822_ _05824_ _05825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_65_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10449__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12590_ memory\[36\]\[15\] memory\[37\]\[15\] _06447_ _06791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13260__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12447__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11541_ _05756_ _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_93_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11810__A2 _06021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14260_ _01299_ clknet_leaf_111_clk_i memory\[15\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13012__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11472_ _05682_ _05685_ _05687_ _05688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09067__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13211_ _05777_ _02604_ _02605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10423_ _05114_ _00255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14191_ _01230_ clknet_leaf_191_clk_i memory\[19\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08814__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13142_ _06844_ _02532_ _02534_ _02536_ _02537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_21_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08152__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10354_ _05014_ memory\[47\]\[4\] _05073_ _05078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12182__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10481__I _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12749__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13073_ memory\[12\]\[22\] memory\[13\]\[22\] _06714_ _02469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10285_ _05032_ _00199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12024_ _06232_ _06233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_168_Right_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_40_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_144_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13079__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_144_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_105_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13975_ _01014_ clknet_leaf_266_clk_i memory\[49\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_105_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11018__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15714_ _00673_ clknet_leaf_315_clk_i memory\[61\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12926_ _06848_ _02323_ _06707_ _02324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_122_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09711__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15645_ _00604_ clknet_leaf_370_clk_i memory\[5\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12857_ _02255_ _02256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_5_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_186_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_16_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11808_ _03120_ _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_51_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12788_ memory\[0\]\[18\] memory\[1\]\[18\] memory\[2\]\[18\] memory\[3\]\[18\] _06709_
+ _06779_ _02188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15576_ _00535_ clknet_leaf_268_clk_i memory\[56\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_154_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14527_ _01566_ clknet_leaf_353_clk_i memory\[24\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11739_ _05951_ _05952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_113_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10860__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14458_ _01497_ clknet_leaf_0_clk_i memory\[21\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13409_ _02337_ _02795_ _02797_ _02799_ _02800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__10592__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14389_ _01428_ clknet_leaf_56_clk_i memory\[1\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_168_3604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11565__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09158__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10612__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08950_ _04214_ memory\[27\]\[15\] _04297_ _04303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_196_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08997__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_138_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07901_ _03714_ _01213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08881_ _04266_ _01641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09230__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_135_Right_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_181_3848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10915__I1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_181_3859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_420_clk_i clknet_5_2__leaf_clk_i clknet_leaf_420_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07832_ _03132_ memory\[7\]\[2\] _03675_ _03678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12312__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07406__S _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07763_ _03641_ _01148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09502_ _04601_ _01927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12111__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07694_ _03129_ memory\[63\]\[1\] _03603_ _03605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09621__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11340__I1 _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_435_clk_i clknet_5_0__leaf_clk_i clknet_leaf_435_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_78_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09433_ _04558_ _01901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10767__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13143__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09364_ _04220_ memory\[33\]\[18\] _04513_ _04522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_192_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08237__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13242__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11479__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12676__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08315_ _03928_ _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_23_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09295_ _04485_ _01836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08246_ _03914_ _01358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09049__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08036__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11598__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12348__A3 _06537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12979__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08177_ _03791_ memory\[29\]\[19\] _03868_ _03878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07128_ _03166_ memory\[13\]\[13\] _03279_ _03283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07059_ _03169_ memory\[16\]\[14\] _03240_ _03245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10007__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10070_ _04912_ _00104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_89_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10906__I1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_102_Right_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09772__I1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07783__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_138_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_398_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13760_ _00799_ clknet_leaf_279_clk_i memory\[14\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10972_ _05018_ memory\[56\]\[6\] _05399_ _05406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12284__A2 _06444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12711_ memory\[48\]\[17\] memory\[49\]\[17\] memory\[50\]\[17\] memory\[51\]\[17\]
+ _06699_ _06839_ _02112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_13691_ _03076_ _00763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10677__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13053__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_100_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15430_ _00389_ clknet_leaf_299_clk_i memory\[52\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12642_ _06831_ _06834_ _06837_ _06841_ _06842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06954__I net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09288__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07051__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15361_ _00320_ clknet_leaf_328_clk_i memory\[50\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12573_ _06411_ _06766_ _06773_ _06774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_136_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14312_ _01351_ clknet_leaf_207_clk_i memory\[17\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11524_ _05736_ _05738_ _05739_ _05740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15292_ _00251_ clknet_leaf_346_clk_i memory\[48\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_110_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1018 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14243_ _01282_ clknet_leaf_279_clk_i memory\[15\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11455_ _03116_ _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11301__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10406_ _05066_ memory\[47\]\[29\] _05095_ _05105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14174_ _01213_ clknet_leaf_350_clk_i memory\[19\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11386_ _05625_ _00707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_110_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13125_ memory\[56\]\[23\] memory\[57\]\[23\] memory\[58\]\[23\] memory\[59\]\[23\]
+ _06827_ _02171_ _02520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_42_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10337_ _05067_ _00216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_163_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13056_ _02170_ _02451_ _02452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09212__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10268_ _05020_ memory\[46\]\[7\] _05006_ _05021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08610__S _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12007_ _05654_ _06211_ _06213_ _06215_ _06216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12132__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10199_ _04595_ memory\[45\]\[10\] _04980_ _04981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07774__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13147__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13958_ _00997_ clknet_leaf_293_clk_i memory\[49\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11322__I1 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09441__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12909_ memory\[56\]\[20\] memory\[57\]\[20\] memory\[58\]\[20\] memory\[59\]\[20\]
+ _06827_ _02171_ _02307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_53_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10587__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13889_ _00928_ clknet_leaf_307_clk_i memory\[11\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15628_ _00587_ clknet_leaf_227_clk_i memory\[58\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11086__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15559_ _00518_ clknet_leaf_233_clk_i memory\[56\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08100_ _03836_ _01290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07896__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09080_ _04208_ memory\[2\]\[12\] _04369_ _04372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_867 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12815__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08031_ _03793_ memory\[12\]\[20\] _03794_ _03795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_135_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09451__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09982_ _04583_ memory\[42\]\[4\] _04861_ _04866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12106__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08933_ _04197_ memory\[27\]\[7\] _04286_ _04294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08520__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09203__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11945__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13138__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11010__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08864_ _04257_ _01633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11710__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07136__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09415__I _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07815_ _03668_ _01173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08795_ _04212_ memory\[25\]\[14\] _04204_ _04213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_84_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_374_clk_i clknet_5_12__leaf_clk_i clknet_leaf_374_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07746_ _03206_ memory\[63\]\[26\] _03625_ _03632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13463__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12897__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11313__I1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07677_ _03595_ _01108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08190__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09416_ _04203_ memory\[34\]\[10\] _04549_ _04550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_176_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_389_clk_i clknet_5_6__leaf_clk_i clknet_leaf_389_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_192_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09347_ _04501_ _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13601__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_117_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09278_ _04476_ _01828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12725__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08229_ _03775_ memory\[17\]\[11\] _03904_ _03906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_312_clk_i clknet_5_11__leaf_clk_i clknet_leaf_312_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_160_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11529__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11121__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11240_ _03317_ memory\[60\]\[4\] _05543_ _05548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10960__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11171_ _05511_ _00606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10122_ _04587_ memory\[44\]\[6\] _04933_ _04940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_327_clk_i clknet_5_10__leaf_clk_i clknet_leaf_327_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09526__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13377__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13048__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10053_ _04903_ _00096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14930_ _01969_ clknet_leaf_72_clk_i memory\[36\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_141_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07046__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07756__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14861_ _01900_ clknet_leaf_51_clk_i memory\[34\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13812_ _00851_ clknet_leaf_115_clk_i memory\[16\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13454__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14792_ _01831_ clknet_leaf_44_clk_i memory\[32\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09261__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13743_ _03103_ _00788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_144_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10955_ _05396_ _00505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13674_ memory\[24\]\[31\] memory\[25\]\[31\] memory\[26\]\[31\] memory\[27\]\[31\]
+ _05742_ _02502_ _03061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10886_ _05359_ _00473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_139_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_139_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15413_ _00372_ clknet_leaf_155_clk_i memory\[51\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12625_ memory\[62\]\[16\] memory\[63\]\[16\] _06557_ _06825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_170_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_14_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10815__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15344_ _00303_ clknet_leaf_146_clk_i memory\[4\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_14_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12556_ _06703_ _06725_ _06741_ _06757_ _06758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_136_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09681__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11507_ _05719_ _05721_ _05722_ _05723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_80_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12487_ memory\[62\]\[14\] memory\[63\]\[14\] _06557_ _06689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15275_ _00234_ clknet_leaf_273_clk_i memory\[47\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14226_ _01265_ clknet_leaf_116_clk_i memory\[12\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11438_ _05653_ _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_151_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11615__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12193__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11966__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14157_ _01196_ clknet_leaf_220_clk_i memory\[7\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11240__I0 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11369_ _03303_ memory\[62\]\[0\] _05616_ _05617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_130_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_69_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13108_ _02501_ _02503_ _02504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_14088_ _01127_ clknet_leaf_223_clk_i memory\[63\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12370__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13039_ memory\[20\]\[21\] memory\[21\]\[21\] _02368_ _02436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_178_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07600_ _03554_ _01072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08580_ _04091_ _01515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_191_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09171__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07531_ _03517_ _01040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13540__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11206__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_176_3758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10110__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07462_ memory\[49\]\[22\] _03355_ _03477_ _03480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13048__I1 net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_176_3769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09201_ _04193_ memory\[31\]\[5\] _04430_ _04436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_493 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11059__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07393_ _03441_ _00978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11759__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09132_ _04399_ _01759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08515__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09063_ _04191_ memory\[2\]\[4\] _04358_ _04363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_346_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08014_ _03171_ _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_5_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09424__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12184__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10780__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11931__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08250__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13359__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13376__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09965_ _04856_ _00055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08916_ _04284_ _01658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07738__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13684__A1 _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09896_ _04633_ memory\[40\]\[28\] _04811_ _04820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08847_ _04247_ memory\[25\]\[31\] _04182_ _04248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08778_ _03152_ _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_58_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07729_ _03181_ memory\[63\]\[18\] _03614_ _03623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08163__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10020__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10740_ _05282_ _00404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_0_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07910__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10671_ memory\[51\]\[25\] _03202_ _05240_ _05246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12098__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12410_ _06603_ _06606_ _06609_ _06613_ _06614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_125_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13390_ memory\[6\]\[27\] memory\[7\]\[27\] _02322_ _02781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_251_clk_i clknet_5_24__leaf_clk_i clknet_leaf_251_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_129_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_11_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11845__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12455__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_97_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12341_ _06545_ _06546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_145_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10754__I _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15060_ _00019_ clknet_leaf_15_clk_i memory\[40\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12272_ memory\[20\]\[10\] memory\[21\]\[10\] _06477_ _06478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_151_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11786__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12175__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14011_ _01050_ clknet_leaf_376_clk_i memory\[59\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11223_ _05538_ _00631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11222__I0 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_75_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_266_clk_i clknet_5_13__leaf_clk_i clknet_leaf_266_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_112_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_70_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11154_ _03367_ memory\[58\]\[28\] _05493_ _05502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12190__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10105_ _04930_ _00121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11085_ _05465_ _00566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07729__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13675__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14913_ _01952_ clknet_leaf_437_clk_i memory\[36\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10036_ _04637_ memory\[42\]\[30\] _04860_ _04894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13506__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14844_ _01883_ clknet_leaf_425_clk_i memory\[34\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07504__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_561 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_204_clk_i clknet_5_30__leaf_clk_i clknet_leaf_204_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_153_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_10__f_clk_i clknet_2_1_0_clk_i clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_81_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_295_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14775_ _01814_ clknet_leaf_86_clk_i memory\[31\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11987_ memory\[24\]\[6\] memory\[25\]\[6\] memory\[26\]\[6\] memory\[27\]\[6\] _05778_
+ _05922_ _06197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08154__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11989__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13726_ _03094_ _00780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10938_ memory\[55\]\[22\] _03193_ _05385_ _05388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12650__A2 _06849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13657_ memory\[38\]\[31\] memory\[39\]\[31\] _05662_ _03044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10865__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10869_ _05052_ memory\[54\]\[22\] _05348_ _05351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12089__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_219_clk_i clknet_5_27__leaf_clk_i clknet_leaf_219_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_128_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12608_ _06607_ _06808_ _06195_ _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_13_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09654__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13588_ memory\[8\]\[30\] memory\[9\]\[30\] memory\[10\]\[30\] memory\[11\]\[30\]
+ _02473_ _05779_ _02976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_171_3666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15327_ _00286_ clknet_leaf_366_clk_i memory\[4\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_30_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12539_ _06445_ _06733_ _06740_ _06741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_121_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15258_ _00217_ clknet_leaf_391_clk_i memory\[46\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14209_ _01248_ clknet_leaf_281_clk_i memory\[12\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15189_ _00148_ clknet_leaf_8_clk_i memory\[44\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08070__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11495__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06962_ net15 _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09750_ _04741_ _02035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13210__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_33_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08701_ _03770_ memory\[24\]\[9\] _04146_ _04156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09681_ _04625_ memory\[37\]\[24\] _04700_ _04705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06893_ _03115_ _03124_ _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_193_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11772__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08632_ _04119_ _01539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12320__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08563_ _04082_ _01507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07514_ _03508_ _01032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08494_ _03768_ memory\[21\]\[8\] _04037_ _04046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07213__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07445_ memory\[49\]\[14\] _03338_ _03466_ _03471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13151__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08245__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07376_ _03432_ _00970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09645__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09115_ _04243_ memory\[2\]\[29\] _04380_ _04390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09046_ _04353_ _01719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_92_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09076__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11904__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_53_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09948_ _04616_ memory\[41\]\[20\] _04847_ _04848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09325__A2 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09879_ _04788_ _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08384__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11910_ memory\[24\]\[5\] memory\[25\]\[5\] memory\[26\]\[5\] memory\[27\]\[5\] _05778_
+ _05922_ _06121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_73_1306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12890_ memory\[24\]\[19\] memory\[25\]\[19\] memory\[26\]\[19\] memory\[27\]\[19\]
+ _06472_ _06611_ _02289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07324__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11841_ memory\[28\]\[4\] memory\[29\]\[4\] _05915_ _06053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_16_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_16_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_17_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14560_ _01599_ clknet_leaf_414_clk_i memory\[25\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11772_ memory\[24\]\[3\] memory\[25\]\[3\] memory\[26\]\[3\] memory\[27\]\[3\] _05778_
+ _05922_ _05985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09884__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13511_ _05724_ _02899_ _02900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10723_ _05273_ _00396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_193_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_190_clk_i clknet_5_29__leaf_clk_i clknet_leaf_190_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14491_ _01530_ clknet_leaf_397_clk_i memory\[22\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06962__I net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13442_ _05700_ _02827_ _02829_ _02831_ _02832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10654_ memory\[51\]\[17\] _03177_ _05229_ _05237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12396__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13373_ memory\[60\]\[27\] memory\[61\]\[27\] _02164_ _02764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_63_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10585_ _05041_ memory\[50\]\[17\] _05192_ _05200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15112_ _00071_ clknet_leaf_29_clk_i memory\[42\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12324_ _06446_ _06524_ _06526_ _06528_ _06529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_161_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12148__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15043_ _00002_ clknet_leaf_433_clk_i memory\[40\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12255_ _05756_ _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13440__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11206_ _03350_ memory\[5\]\[20\] _05529_ _05530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_107_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12186_ _05731_ _06385_ _06392_ _06393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_11137_ _05470_ _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_78_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11068_ _05456_ _00558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08375__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13236__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10019_ _04885_ _00080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12140__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_143_clk_i clknet_5_19__leaf_clk_i clknet_leaf_143_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10182__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14827_ _01866_ clknet_leaf_45_clk_i memory\[33\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14758_ _01797_ clknet_leaf_132_clk_i memory\[31\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09875__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13709_ _03085_ _00772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_158_clk_i clknet_5_24__leaf_clk_i clknet_leaf_158_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14689_ _01728_ clknet_leaf_359_clk_i memory\[2\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07968__I _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07230_ _03347_ _00909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09627__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11809__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07161_ _03215_ memory\[13\]\[29\] _03290_ _03300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07092_ _03218_ memory\[16\]\[30\] _03228_ _03262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12139__A1 _06292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_188_3982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_188_3993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09802_ _04769_ _02059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12114__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13639__A1 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07994_ _03769_ _01251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06945_ _03164_ _00807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09733_ _04732_ _02027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09664_ _04608_ memory\[37\]\[16\] _04689_ _04696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_2_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08615_ memory\[23\]\[0\] _03303_ _04110_ _04111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12985__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09595_ _04659_ _01962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08118__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08039__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08546_ _03746_ memory\[22\]\[0\] _04073_ _04074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08669__I1 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08477_ _04036_ _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_175_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07428_ memory\[49\]\[6\] _03321_ _03455_ _03462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_46_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_162_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11425__I0 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07359_ _03423_ _00962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_94_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_116_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_149_Right_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10370_ _05086_ _00230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_60_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_243_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12733__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09029_ _04224_ memory\[28\]\[20\] _04344_ _04345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13422__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12040_ memory\[46\]\[7\] memory\[47\]\[7\] _05907_ _06249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_60_clk_i clknet_5_17__leaf_clk_i clknet_leaf_60_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13991_ _01030_ clknet_leaf_296_clk_i memory\[59\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12302__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15730_ _00689_ clknet_leaf_146_clk_i memory\[61\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12942_ _02339_ _02340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10164__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15661_ _00620_ clknet_leaf_252_clk_i memory\[5\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12895__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12873_ memory\[38\]\[19\] memory\[39\]\[19\] _06728_ _02272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_75_clk_i clknet_5_17__leaf_clk_i clknet_leaf_75_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14612_ _01651_ clknet_leaf_95_clk_i memory\[26\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11824_ _05699_ _06023_ _06035_ _06036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_15592_ _00551_ clknet_leaf_232_clk_i memory\[57\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_103_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_190_4028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12908__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12161__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10616__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14543_ _01582_ clknet_leaf_185_clk_i memory\[24\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11755_ memory\[38\]\[3\] memory\[39\]\[3\] _05737_ _05968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_83_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_83_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07332__I1 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10706_ _05264_ _00388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_193_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14474_ _01513_ clknet_leaf_197_clk_i memory\[22\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09609__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11686_ memory\[38\]\[2\] memory\[39\]\[2\] _05737_ _05900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13425_ memory\[20\]\[27\] memory\[21\]\[27\] _02368_ _02816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10637_ memory\[51\]\[9\] _03152_ _05218_ _05228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09709__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13356_ _02747_ _02748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10568_ _05024_ memory\[50\]\[9\] _05181_ _05191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_116_Right_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_13_clk_i clknet_5_5__leaf_clk_i clknet_leaf_13_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12307_ memory\[0\]\[11\] memory\[1\]\[11\] memory\[2\]\[11\] memory\[3\]\[11\] _06020_
+ _06090_ _06512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_84_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10499_ _05154_ _00291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13287_ _02213_ _02679_ _02352_ _02680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_121_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15026_ _02065_ clknet_leaf_56_clk_i memory\[3\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12238_ _06428_ _06436_ _06443_ _06444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08596__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11974__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_166_3565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12169_ _06031_ _06375_ _06376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
Xclkbuf_leaf_28_clk_i clknet_5_6__leaf_clk_i clknet_leaf_28_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_183_3890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_445_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08348__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11727__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 address_i[4] net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_56_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_155_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08400_ _03810_ memory\[1\]\[28\] _03987_ _03996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09380_ _04530_ _01876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_192_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09848__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_135_Left_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08331_ _03959_ _01398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08520__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_145_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11214__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08262_ _03808_ memory\[17\]\[27\] _03915_ _03923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07213_ _03165_ _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_160_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08193_ _03886_ _01333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07144_ _03291_ _00879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_5_23__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09619__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_41_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07075_ _03253_ _00848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_144_Left_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_65_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13324__A3 _02715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_7_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10394__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input37_I data_i[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07977_ _03134_ _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09716_ _04723_ _02019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_06928_ _03151_ _00803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_87_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09647_ _04591_ memory\[37\]\[8\] _04678_ _04687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_Left_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_48_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_48_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09578_ _04650_ _01954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_65_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_77_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08529_ _04064_ _01491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08511__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11540_ _03112_ _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11471_ _05686_ _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09067__I1 memory\[2\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07078__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13210_ memory\[8\]\[24\] memory\[9\]\[24\] memory\[10\]\[24\] memory\[11\]\[24\]
+ _02473_ _05779_ _02604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_150_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10422_ _05014_ memory\[48\]\[4\] _05109_ _05114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09529__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08433__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14190_ _01229_ clknet_leaf_196_clk_i memory\[19\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_394_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_162_Left_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13141_ _06851_ _02535_ _02536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10621__I1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10353_ _05077_ _00222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13072_ _06844_ _02463_ _02465_ _02467_ _02468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_103_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10284_ _05031_ memory\[46\]\[12\] _05027_ _05032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12523__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11794__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12023_ memory\[12\]\[7\] memory\[13\]\[7\] _06025_ _06232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10385__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_144_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11807__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_144_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11709__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10137__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13974_ _01013_ clknet_leaf_263_clk_i memory\[49\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_105_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_171_Left_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_161_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15713_ _00672_ clknet_leaf_323_clk_i memory\[61\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12925_ memory\[6\]\[20\] memory\[7\]\[20\] _02322_ _02323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13514__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15644_ _00603_ clknet_leaf_370_clk_i memory\[5\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12856_ memory\[4\]\[19\] memory\[5\]\[19\] _06845_ _02255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08608__S _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11542__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11807_ _05705_ _06017_ _06018_ _06019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15575_ _00534_ clknet_leaf_253_clk_i memory\[56\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12787_ _06848_ _02186_ _06707_ _02187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_111_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07305__I1 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11034__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14526_ _01565_ clknet_leaf_353_clk_i memory\[24\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11738_ memory\[4\]\[3\] memory\[5\]\[3\] _05702_ _05951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14457_ _01496_ clknet_leaf_98_clk_i memory\[21\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10873__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11669_ _05882_ _05883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XPHY_EDGE_ROW_180_Left_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07069__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13408_ _02344_ _02798_ _02799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_114_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09439__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13469__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14388_ _01427_ clknet_leaf_57_clk_i memory\[1\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_4_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13339_ _02319_ _02723_ _02730_ _02731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_84_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_139_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_3930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_122_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13306__A3 _02698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_185_3941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08569__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15009_ _02048_ clknet_leaf_340_clk_i memory\[3\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07900_ _03132_ memory\[19\]\[2\] _03711_ _03714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08880_ _04212_ memory\[26\]\[14\] _04261_ _04266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_181_3849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07831_ _03677_ _01180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10128__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07762_ _03129_ memory\[6\]\[1\] _03639_ _03641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09902__S _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09501_ _04600_ memory\[35\]\[12\] _04596_ _04601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07693_ _03604_ _01115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10679__I1 _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08741__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07544__I1 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09432_ _04220_ memory\[34\]\[18\] _04549_ _04558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_52_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09363_ _04521_ _01868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12676__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08314_ _03950_ _01390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_19_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_23_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09294_ _04218_ memory\[32\]\[17\] _04477_ _04485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08245_ _03791_ memory\[17\]\[19\] _03904_ _03914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08176_ _03877_ _01325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_162_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12348__A4 _06552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07127_ _03282_ _00871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07058_ _03244_ _00840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10367__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_89_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09084__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07232__I0 memory\[39\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11119__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09812__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10971_ _05405_ _00512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12284__A3 _06466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13334__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12710_ _06835_ _02110_ _06287_ _02111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_35_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08428__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13690_ _03303_ memory\[9\]\[0\] _03075_ _03076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07332__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_100_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12641_ _06838_ _06840_ _06841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_182_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_80_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15360_ _00319_ clknet_leaf_329_clk_i memory\[50\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12572_ _06142_ _06768_ _06770_ _06772_ _06773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_108_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14311_ _01350_ clknet_leaf_205_clk_i memory\[17\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12992__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11523_ _05686_ _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10693__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15291_ _00250_ clknet_leaf_392_clk_i memory\[47\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09259__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06970__I net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14242_ _01281_ clknet_leaf_281_clk_i memory\[15\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08163__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11454_ _05669_ _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_85_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12744__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10405_ _05104_ _00247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14173_ _01212_ clknet_leaf_363_clk_i memory\[19\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11385_ _03325_ memory\[62\]\[8\] _05616_ _05625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_104_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_140_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13124_ _02167_ _02518_ _06690_ _02519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_81_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10336_ _05066_ memory\[46\]\[29\] _05048_ _05067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12413__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13055_ memory\[56\]\[22\] memory\[57\]\[22\] memory\[58\]\[22\] memory\[59\]\[22\]
+ _06827_ _02171_ _02451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10267_ _03146_ _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_163_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10358__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12006_ _05668_ _06214_ _06215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07223__I0 memory\[39\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07507__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10198_ _04968_ _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_84_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08971__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09722__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13957_ _00996_ clknet_leaf_317_clk_i memory\[49\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12908_ _02167_ _02305_ _06690_ _02306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_159_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10530__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08338__S _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13888_ _00927_ clknet_leaf_307_clk_i memory\[11\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12107__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09521__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07242__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15627_ _00586_ clknet_leaf_230_clk_i memory\[58\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_65_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12839_ _02238_ net49 _06491_ _02239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08137__I _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15558_ _00517_ clknet_leaf_229_clk_i memory\[56\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14509_ _01548_ clknet_leaf_174_clk_i memory\[23\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12983__A1 _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15489_ _00448_ clknet_leaf_328_clk_i memory\[54\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08030_ _03751_ _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_126_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09169__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06880__I net4 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput30 data_i[30] net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_4_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09981_ _04865_ _00062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08932_ _04293_ _01665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07214__I0 memory\[39\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12594__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08863_ _04195_ memory\[26\]\[6\] _04250_ _04257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_36_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07814_ _03206_ memory\[6\]\[26\] _03661_ _03668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_342_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08794_ _03168_ _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07216__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_84_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07745_ _03631_ _01140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10778__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08714__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07517__I1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12897__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08248__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07676_ _03203_ memory\[10\]\[25\] _03589_ _03595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10521__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09415_ _04537_ _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_62_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09346_ _04512_ _01860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_1300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09277_ _04201_ memory\[32\]\[9\] _04466_ _04476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11402__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_99_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08228_ _03905_ _01349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08159_ _03772_ memory\[29\]\[10\] _03868_ _03869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10018__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09807__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11170_ _03315_ memory\[5\]\[3\] _05507_ _05511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10121_ _04939_ _00128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12233__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_output68_I net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07205__I0 memory\[39\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10052_ _04585_ memory\[43\]\[5\] _04897_ _04903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14860_ _01899_ clknet_leaf_51_clk_i memory\[34\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12337__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13811_ _00850_ clknet_leaf_117_clk_i memory\[16\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13572__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14791_ _01830_ clknet_leaf_50_clk_i memory\[32\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13742_ _03361_ memory\[9\]\[25\] _03097_ _03103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10954_ memory\[55\]\[30\] _03217_ _05362_ _05396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13673_ _02498_ _03059_ _05665_ _03060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_183_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_168_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10885_ _05068_ memory\[54\]\[30\] _05325_ _05359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15412_ _00371_ clknet_leaf_155_clk_i memory\[51\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A1 _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12624_ _06823_ _06824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12916__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_14_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15343_ _00302_ clknet_leaf_254_clk_i memory\[4\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12555_ _06467_ _06748_ _06756_ _06757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_93_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_0_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_123_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11506_ _05664_ _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_117_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07692__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15274_ _00233_ clknet_leaf_275_clk_i memory\[47\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_41_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12486_ _06687_ _06688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_184_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14225_ _01264_ clknet_leaf_118_clk_i memory\[12\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11437_ _05652_ _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_34_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10579__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09717__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14156_ _01195_ clknet_leaf_220_clk_i memory\[7\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_434_clk_i clknet_5_0__leaf_clk_i clknet_leaf_434_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08621__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11368_ _05615_ _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_120_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13107_ memory\[24\]\[22\] memory\[25\]\[22\] memory\[26\]\[22\] memory\[27\]\[22\]
+ _02363_ _02502_ _02503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_130_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10319_ _05055_ _00210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14087_ _01126_ clknet_leaf_228_clk_i memory\[63\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11299_ _05578_ _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13142__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09197__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13038_ _06603_ _02430_ _02432_ _02434_ _02435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08944__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10751__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10598__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14989_ _02028_ clknet_leaf_43_clk_i memory\[38\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_18_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07530_ memory\[59\]\[21\] _03353_ _03515_ _03517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08068__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10503__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07461_ _03479_ _01008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_176_3759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09200_ _04435_ _01791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13702__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06883__A1 _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07392_ _03197_ memory\[8\]\[23\] _03437_ _03441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07700__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09131_ _04191_ memory\[30\]\[4\] _04394_ _04399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12318__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11222__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09062_ _04362_ _01726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_60_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08013_ _03782_ _01257_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12117__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_12_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09627__S _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12053__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09964_ _04633_ memory\[41\]\[28\] _04847_ _04856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07147__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13133__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08915_ _04247_ memory\[26\]\[31\] _04249_ _04284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09895_ _04819_ _00022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08935__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11695__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08846_ _03220_ _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_100_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_51_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09362__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08777_ _04200_ _01603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07728_ _03622_ _01132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09360__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07659_ _03178_ memory\[10\]\[17\] _03578_ _03586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_137_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10670_ _05245_ _00371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08706__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09329_ _04185_ memory\[33\]\[1\] _04502_ _04504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12340_ memory\[20\]\[11\] memory\[21\]\[11\] _06477_ _06545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07674__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12271_ _05784_ _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_151_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14010_ _01049_ clknet_leaf_380_clk_i memory\[59\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_75_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_107_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11222_ _03367_ memory\[5\]\[28\] _05529_ _05538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08441__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_13_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11153_ _05501_ _00598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10981__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07057__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13124__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09179__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10104_ _04637_ memory\[43\]\[30\] _04896_ _04930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11084_ _05062_ memory\[57\]\[27\] _05457_ _05465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14912_ _01951_ clknet_leaf_424_clk_i memory\[36\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10035_ _04893_ _00088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10733__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14843_ _01882_ clknet_leaf_0_clk_i memory\[33\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11307__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_238_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10211__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14774_ _01813_ clknet_leaf_86_clk_i memory\[31\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11986_ _05918_ _06194_ _06195_ _06196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_187_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13725_ _03344_ memory\[9\]\[17\] _03086_ _03094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10937_ _05387_ _00496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13656_ _03042_ _03043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10868_ _05350_ _00464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09103__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12607_ memory\[30\]\[15\] memory\[31\]\[15\] _06193_ _06808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_155_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13587_ _05772_ _02974_ _05775_ _02975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11042__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10799_ _05050_ memory\[53\]\[21\] _05312_ _05314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15326_ _00285_ clknet_leaf_339_clk_i memory\[4\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11610__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12538_ _06318_ _06735_ _06737_ _06739_ _06740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_14_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13738__I0 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_112_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10881__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15257_ _00216_ clknet_leaf_385_clk_i memory\[46\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12469_ memory\[30\]\[13\] memory\[31\]\[13\] _06193_ _06672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_373_clk_i clknet_5_12__leaf_clk_i clknet_leaf_373_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14208_ _01247_ clknet_leaf_279_clk_i memory\[12\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09447__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12797__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15188_ _00147_ clknet_leaf_15_clk_i memory\[44\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14139_ _01178_ clknet_leaf_393_clk_i memory\[6\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10972__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13115__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06961_ _03176_ _00811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_388_clk_i clknet_5_6__leaf_clk_i clknet_leaf_388_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13210__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08700_ _04155_ _01571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09680_ _04704_ _02002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06892_ _03118_ _03123_ _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__10724__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09590__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11772__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08631_ memory\[23\]\[8\] _03325_ _04110_ _04119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_311_clk_i clknet_5_11__leaf_clk_i clknet_leaf_311_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12400__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08562_ _03768_ memory\[22\]\[8\] _04073_ _04082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09910__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07513_ memory\[59\]\[13\] _03336_ _03504_ _03508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_18_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08493_ _04045_ _01474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07444_ _03470_ _01000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_186_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08526__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_326_clk_i clknet_5_10__leaf_clk_i clknet_leaf_326_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12929__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07430__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07375_ _03172_ memory\[8\]\[15\] _03426_ _03432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12048__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09114_ _04389_ _01751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11601__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13729__I0 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09045_ _04241_ memory\[28\]\[28\] _04344_ _04353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_57_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07408__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13354__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12788__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_92_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12291__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_187_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_53_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_53_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08060__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09947_ _04824_ _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_70_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13607__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09878_ _04810_ _00014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09092__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07605__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08829_ _04235_ memory\[25\]\[25\] _04225_ _04236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13409__A2 _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11127__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11840_ _05731_ _06044_ _06051_ _06052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_135_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09333__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_16_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_36_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11771_ _05918_ _05983_ _05775_ _05984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10966__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11140__I0 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13342__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13510_ memory\[48\]\[29\] memory\[49\]\[29\] memory\[50\]\[29\] memory\[51\]\[29\]
+ _05725_ _05726_ _02899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10722_ _05041_ memory\[52\]\[17\] _05265_ _05273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_192_4070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11840__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14490_ _01529_ clknet_leaf_398_clk_i memory\[22\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07340__S _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13441_ _05710_ _02830_ _02831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_193_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10653_ _05236_ _00363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_153_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07647__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13372_ _02763_ _00757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10584_ _05199_ _00331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_106_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15111_ _00070_ clknet_leaf_22_clk_i memory\[42\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12323_ _06453_ _06527_ _06528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_106_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Left_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_106_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09267__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15042_ _00001_ clknet_leaf_433_clk_i memory\[40\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08171__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12254_ memory\[46\]\[10\] memory\[47\]\[10\] _05907_ _06460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13440__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07024__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11205_ _05506_ _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08072__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12185_ _06318_ _06387_ _06389_ _06391_ _06392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_120_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11136_ _05492_ _00590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11659__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11067_ _05045_ memory\[57\]\[19\] _05446_ _05456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07515__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10018_ _04619_ memory\[42\]\[21\] _04883_ _04885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_48_Left_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_389_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14826_ _01865_ clknet_leaf_44_clk_i memory\[33\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_125_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_125_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09730__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14757_ _01796_ clknet_leaf_404_clk_i memory\[31\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12084__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11131__I0 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11969_ memory\[32\]\[6\] memory\[33\]\[6\] memory\[34\]\[6\] memory\[35\]\[6\] _05742_
+ _05743_ _06179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_153_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_3707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13708_ _03327_ memory\[9\]\[9\] _03075_ _03085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07886__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11831__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14688_ _01727_ clknet_leaf_359_clk_i memory\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08346__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13639_ _03450_ _03018_ _03025_ _03026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_172_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_441_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07160_ _03299_ _00887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07638__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_13__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_57_Left_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15309_ _00268_ clknet_leaf_257_clk_i memory\[48\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_171_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07091_ _03261_ _00856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09177__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10116__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09801_ memory\[3\]\[16\] _03174_ _04762_ _04769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_1_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07810__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07993_ _03768_ memory\[12\]\[8\] _03752_ _03769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13427__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09732_ _04608_ memory\[38\]\[16\] _04725_ _04732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13195__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06944_ _03163_ memory\[14\]\[12\] _03157_ _03164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_250_clk_i clknet_5_25__leaf_clk_i clknet_leaf_250_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09563__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_66_Left_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09663_ _04695_ _01994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_2_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_2_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08614_ _04109_ _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_96_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09594_ _04606_ memory\[36\]\[15\] _04653_ _04659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09315__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08545_ _04072_ _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12075__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10786__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11822__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08256__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08476_ _03225_ _03266_ _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_148_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07427_ _03461_ _00992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_92_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_45_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13575__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07358_ _03147_ memory\[8\]\[7\] _03415_ _03423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_94_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07289_ _03386_ _00929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_115_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09028_ _04321_ _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11189__I0 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_203_clk_i clknet_5_30__leaf_clk_i clknet_leaf_203_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_143_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13422__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11889__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10026__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_9_clk_i clknet_5_5__leaf_clk_i clknet_leaf_9_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
Xclkbuf_leaf_218_clk_i clknet_5_27__leaf_clk_i clknet_leaf_218_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13990_ _01029_ clknet_leaf_236_clk_i memory\[59\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_output50_I net50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_146_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12941_ memory\[36\]\[20\] memory\[37\]\[20\] _02338_ _02339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_390_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15660_ _00619_ clknet_leaf_252_clk_i memory\[5\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12872_ _02270_ _02271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__09550__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14611_ _01650_ clknet_leaf_96_clk_i memory\[26\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13580__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11823_ _06024_ _06027_ _06030_ _06034_ _06035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12975__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15591_ _00550_ clknet_leaf_233_clk_i memory\[57\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_190_4029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14542_ _01581_ clknet_leaf_185_clk_i memory\[24\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12161__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11754_ _05966_ _05967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10616__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_83_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10705_ _05024_ memory\[52\]\[9\] _05254_ _05264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14473_ _01512_ clknet_leaf_175_clk_i memory\[22\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11685_ _05898_ _05899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_13424_ _02494_ _02810_ _02812_ _02814_ _02815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_37_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10636_ _05227_ _00355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13355_ memory\[28\]\[26\] memory\[29\]\[26\] _02495_ _02747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11672__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10567_ _05190_ _00323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12306_ _06159_ _06510_ _06018_ _06511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13286_ memory\[46\]\[25\] memory\[47\]\[25\] _02487_ _02679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10498_ _05022_ memory\[4\]\[8\] _05145_ _05154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15025_ _02064_ clknet_leaf_89_clk_i memory\[3\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12237_ _06024_ _06438_ _06440_ _06442_ _06443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__12215__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_166_3566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12168_ memory\[8\]\[9\] memory\[9\]\[9\] memory\[10\]\[9\] memory\[11\]\[9\] _05893_
+ _06032_ _06375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_120_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13247__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13177__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11119_ _03332_ memory\[58\]\[11\] _05482_ _05484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_183_3891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12151__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12099_ _06031_ _06306_ _06307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_127_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_127_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09524__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07245__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11727__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 address_i[5] net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_127_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11990__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_118_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14809_ _01848_ clknet_leaf_69_clk_i memory\[32\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_135_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11104__I0 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15789_ _00748_ clknet_leaf_260_clk_i net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08330_ _03808_ memory\[18\]\[27\] _03951_ _03959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07859__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08076__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08261_ _03922_ _01365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13557__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07212_ _03335_ _00903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08804__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08192_ _03806_ memory\[29\]\[26\] _03879_ _03886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07143_ _03187_ memory\[13\]\[20\] _03290_ _03291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08284__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_41_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07074_ _03191_ memory\[16\]\[21\] _03251_ _03253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07219__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09635__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_58_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_22_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13665__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07976_ _03757_ _01245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07155__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09715_ _04591_ memory\[38\]\[8\] _04714_ _04723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06927_ _03150_ memory\[14\]\[8\] _03126_ _03151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12996__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_87_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09646_ _04686_ _01986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_48_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_182_Right_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12795__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09577_ _04589_ memory\[36\]\[7\] _04642_ _04650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08528_ _03802_ memory\[21\]\[24\] _04059_ _04064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08459_ _04027_ _01458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_14_Right_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_80_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11470_ _03113_ _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_92_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08714__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10421_ _05113_ _00254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_337_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12220__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11140__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_142_clk_i clknet_5_19__leaf_clk_i clknet_leaf_142_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13140_ memory\[0\]\[23\] memory\[1\]\[23\] memory\[2\]\[23\] memory\[3\]\[23\] _06709_
+ _06779_ _02535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_60_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10352_ _05012_ memory\[47\]\[3\] _05073_ _05077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08027__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13071_ _06851_ _02466_ _02467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_104_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10283_ _03162_ _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_148_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12022_ _06155_ _06226_ _06228_ _06230_ _06231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_40_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_23_Right_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_157_clk_i clknet_5_24__leaf_clk_i clknet_leaf_157_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_144_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07065__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11709__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13973_ _01012_ clknet_leaf_264_clk_i memory\[49\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_161_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12924_ _05661_ _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15712_ _00671_ clknet_leaf_323_clk_i memory\[61\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09280__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15643_ _00602_ clknet_leaf_376_clk_i memory\[58\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12855_ _06411_ _02246_ _02253_ _02254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_38_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11315__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11806_ _05686_ _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_84_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15574_ _00533_ clknet_leaf_159_clk_i memory\[56\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12786_ memory\[6\]\[18\] memory\[7\]\[18\] _06431_ _02186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_32_Right_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14525_ _01564_ clknet_leaf_407_clk_i memory\[24\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_113_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11737_ _05651_ _05942_ _05949_ _05950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_25_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_3_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13539__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14456_ _01495_ clknet_leaf_92_clk_i memory\[21\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11668_ memory\[4\]\[2\] memory\[5\]\[2\] _05702_ _05882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_153_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13407_ memory\[32\]\[27\] memory\[33\]\[27\] memory\[34\]\[27\] memory\[35\]\[27\]
+ _02205_ _02345_ _02798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08266__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10619_ memory\[51\]\[0\] _03110_ _05218_ _05219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12211__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14387_ _01426_ clknet_leaf_139_clk_i memory\[1\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12062__I1 net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11645__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11599_ _05682_ _05813_ _05687_ _05814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_98_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10073__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13338_ _05768_ _02725_ _02727_ _02729_ _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_3_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08018__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13269_ memory\[12\]\[25\] memory\[13\]\[25\] _05769_ _02662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_185_3942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_41_Right_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_62_1350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15008_ _02047_ clknet_leaf_341_clk_i memory\[3\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09455__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_61_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07830_ _03129_ memory\[7\]\[1\] _03675_ _03677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_159_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07761_ _03640_ _01147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09500_ _03162_ _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07692_ _03111_ memory\[63\]\[0\] _03603_ _03604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09431_ _04557_ _01900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11733__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_286_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_50_Right_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09362_ _04218_ memory\[33\]\[17\] _04513_ _04521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08313_ _03791_ memory\[18\]\[19\] _03940_ _03950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_19_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12450__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09293_ _04484_ _01835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08244_ _03913_ _01357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08534__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_60_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08175_ _03789_ memory\[29\]\[18\] _03868_ _03877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07126_ _03163_ memory\[13\]\[12\] _03279_ _03282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08009__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07057_ _03166_ memory\[16\]\[13\] _03240_ _03244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_74_clk_i clknet_5_16__leaf_clk_i clknet_leaf_74_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_113_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06989__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07480__I1 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09757__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_89_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07232__I1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09164__I _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12269__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_89_clk_i clknet_5_20__leaf_clk_i clknet_leaf_89_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07959_ _03744_ _01241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_925 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_74_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10970_ _05016_ memory\[56\]\[5\] _05399_ _05405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_97_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07613__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12284__A4 _06489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09629_ net76 _03305_ _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_74_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_clk_i clknet_5_16__leaf_clk_i clknet_leaf_12_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11135__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_100_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12640_ memory\[48\]\[16\] memory\[49\]\[16\] memory\[50\]\[16\] memory\[51\]\[16\]
+ _06699_ _06839_ _06840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_155_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_80_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07299__I1 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08496__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12571_ _06149_ _06771_ _06772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_66_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14310_ _01349_ clknet_leaf_205_clk_i memory\[17\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11522_ memory\[38\]\[0\] memory\[39\]\[0\] _05737_ _05738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15290_ _00249_ clknet_leaf_392_clk_i memory\[47\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_27_clk_i clknet_5_4__leaf_clk_i clknet_leaf_27_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_109_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_191_882 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14241_ _01280_ clknet_leaf_280_clk_i memory\[15\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_190_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08248__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11453_ _03119_ _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_12
XFILLER_0_68_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10404_ _05064_ memory\[47\]\[28\] _05095_ _05104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14172_ _01211_ clknet_leaf_367_clk_i memory\[19\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11384_ _05624_ _00706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13123_ memory\[62\]\[23\] memory\[63\]\[23\] _02448_ _02518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_78_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10335_ _03214_ _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_115_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06899__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09275__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13054_ _02167_ _02449_ _06690_ _02450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10266_ _05019_ _00193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11818__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12005_ memory\[56\]\[7\] memory\[57\]\[7\] memory\[58\]\[7\] memory\[59\]\[7\] _06138_
+ _05671_ _06214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__07223__I1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08420__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10197_ _04979_ _00164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11858__I1 net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08619__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13956_ _00995_ clknet_leaf_317_clk_i memory\[49\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07523__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09920__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12907_ memory\[62\]\[20\] memory\[63\]\[20\] _06557_ _02305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13887_ _00926_ clknet_leaf_311_clk_i memory\[11\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_75_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12107__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15626_ _00585_ clknet_leaf_230_clk_i memory\[58\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12838_ _02183_ _02200_ _02221_ _02237_ _02238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_185_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_186_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12432__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12769_ _02167_ _02168_ _06690_ _02169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15557_ _00516_ clknet_leaf_319_clk_i memory\[56\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_189_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_71_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14508_ _01547_ clknet_leaf_174_clk_i memory\[23\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12983__A2 _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_126_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15488_ _00447_ clknet_leaf_333_clk_i memory\[54\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_16_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08354__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08239__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput20 data_i[21] net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14439_ _01478_ clknet_leaf_189_clk_i memory\[21\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput31 data_i[31] net31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10046__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_1__f_clk_i clknet_2_0_0_clk_i clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09980_ _04581_ memory\[42\]\[3\] _04861_ _04865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07462__I1 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07992__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09185__S _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08931_ _04195_ memory\[27\]\[6\] _04286_ _04293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12499__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12403__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08862_ _04256_ _01632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07214__I1 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12594__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07813_ _03667_ _01172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08793_ _04211_ _01608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07744_ _03203_ memory\[63\]\[25\] _03625_ _03631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07675_ _03594_ _01107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09414_ _04548_ _01892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09345_ _04201_ memory\[33\]\[9\] _04502_ _04512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08478__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10794__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_34_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08264__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09276_ _04475_ _01827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08227_ _03772_ memory\[17\]\[10\] _03904_ _03905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09978__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_880 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08158_ _03856_ _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08063__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07109_ _03138_ memory\[13\]\[4\] _03268_ _03273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08089_ _03772_ memory\[15\]\[10\] _03830_ _03831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07453__I1 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_101_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10120_ _04585_ memory\[44\]\[5\] _04933_ _04939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08402__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10051_ _04902_ _00095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10034__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07205__I1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_73_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11162__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06964__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13810_ _00849_ clknet_leaf_102_clk_i memory\[16\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12337__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14790_ _01829_ clknet_leaf_46_clk_i memory\[32\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08439__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_11_Left_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09902__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13741_ _03102_ _00787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12662__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10953_ _05395_ _00504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13672_ memory\[30\]\[31\] memory\[31\]\[31\] _05737_ _03059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_167_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10884_ _05358_ _00472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07142__I _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_139_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12623_ memory\[60\]\[16\] memory\[61\]\[16\] _06273_ _06823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15411_ _00370_ clknet_leaf_153_clk_i memory\[51\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12414__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06892__A2 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15342_ _00301_ clknet_leaf_252_clk_i memory\[4\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12554_ _06476_ _06750_ _06753_ _06755_ _06756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_156_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11505_ memory\[14\]\[0\] memory\[15\]\[0\] _05720_ _05721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15273_ _00232_ clknet_leaf_277_clk_i memory\[47\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_117_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10209__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12485_ memory\[60\]\[14\] memory\[61\]\[14\] _06273_ _06687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_117_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_20_Left_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_151_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10028__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14224_ _01263_ clknet_leaf_116_clk_i memory\[12\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11436_ _03116_ _03264_ _05652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_0_110_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_234_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14155_ _01194_ clknet_leaf_221_clk_i memory\[7\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12424__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11367_ _03124_ _03490_ _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_123_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13106_ _03747_ _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10318_ _05054_ memory\[46\]\[23\] _05048_ _05055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_130_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14086_ _01125_ clknet_leaf_222_clk_i memory\[63\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11298_ _03266_ _03490_ _05578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13037_ _06610_ _02433_ _02434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10249_ _03128_ _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07317__I _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10879__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13525__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14988_ _02027_ clknet_leaf_43_clk_i memory\[38\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13939_ _00978_ clknet_leaf_123_clk_i memory\[8\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12653__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07460_ memory\[49\]\[21\] _03353_ _03477_ _03479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12405__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15609_ _00568_ clknet_leaf_270_clk_i memory\[57\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07391_ _03440_ _00977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06883__A2 _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09130_ _04398_ _01758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_57_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08084__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07132__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_893 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09061_ _04189_ memory\[2\]\[3\] _04358_ _04362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08880__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08012_ _03781_ memory\[12\]\[14\] _03773_ _03782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09908__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_38_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07428__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11458__B _05666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_4_Right_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09963_ _04855_ _00054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08914_ _04283_ _01657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09894_ _04631_ memory\[40\]\[27\] _04811_ _04819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09643__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13673__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08845_ _04246_ _01625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12892__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_436_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_51_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08776_ _04199_ memory\[25\]\[8\] _04183_ _04200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input12_I data_i[14] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07163__S _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07727_ _03178_ memory\[63\]\[17\] _03614_ _03622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_2__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08699__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13692__I0 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07658_ _03585_ _01099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11998__A3 _06190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_183_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07371__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07589_ _03548_ _01067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11413__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09328_ _04503_ _01851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10958__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_69_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09259_ _04181_ memory\[32\]\[0\] _04466_ _04467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09818__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12270_ _05747_ _06476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__08722__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11221_ _05537_ _00630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07426__I1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_75_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10430__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07338__S _03378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11152_ _03365_ memory\[58\]\[27\] _05493_ _05501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10103_ _04929_ _00120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11083_ _05464_ _00565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09553__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14911_ _01950_ clknet_leaf_436_clk_i memory\[36\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10034_ _04635_ memory\[42\]\[29\] _04883_ _04893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12978__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10699__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12883__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13075__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06976__I _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14842_ _01881_ clknet_leaf_5_clk_i memory\[33\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08169__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11985_ _05664_ _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14773_ _01812_ clknet_leaf_87_clk_i memory\[31\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_158_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13724_ _03093_ _00779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_158_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10936_ memory\[55\]\[21\] _03190_ _05385_ _05387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07362__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13655_ memory\[36\]\[31\] memory\[37\]\[31\] _05656_ _03042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10867_ _05050_ memory\[54\]\[21\] _05348_ _05350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12606_ _06806_ _06807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13586_ memory\[14\]\[30\] memory\[15\]\[30\] _05773_ _02974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10798_ _05313_ _00431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15325_ _00284_ clknet_leaf_341_clk_i memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12537_ _06325_ _06738_ _06739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_30_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09728__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12468_ _06670_ _06671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_132_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15256_ _00215_ clknet_leaf_39_clk_i memory\[46\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_385_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11419_ _03359_ memory\[62\]\[24\] _05638_ _05643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14207_ _01246_ clknet_leaf_374_clk_i memory\[12\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12797__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15187_ _00146_ clknet_leaf_14_clk_i memory\[44\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12399_ _05653_ _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__07248__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14138_ _01177_ clknet_leaf_393_clk_i memory\[6\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14069_ _01108_ clknet_leaf_113_clk_i memory\[10\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06960_ _03175_ memory\[14\]\[16\] _03157_ _03176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input4_I address_i[3] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06891_ _03121_ _03122_ _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__12874__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08630_ _04118_ _01538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10402__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08561_ _04081_ _01506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12626__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13713__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10488__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07512_ _03507_ _01031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08492_ _03766_ memory\[21\]\[7\] _04037_ _04045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_18_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08807__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11741__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07443_ memory\[49\]\[13\] _03336_ _03466_ _03470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_175_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07374_ _03431_ _00969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07105__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_190_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_130_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09113_ _04241_ memory\[2\]\[28\] _04380_ _04389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08853__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09044_ _04352_ _01718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13668__B _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08542__S _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11967__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12788__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_92_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_92_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08341__I _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06997__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09946_ _04846_ _00046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_70_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09373__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11916__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06919__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09877_ _04614_ memory\[40\]\[19\] _04800_ _04810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11408__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10312__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08828_ _03202_ _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07592__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_79_Right_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08759_ _04188_ _01597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13623__S _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11770_ memory\[30\]\[3\] memory\[31\]\[3\] _05773_ _05983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07344__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13290__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_433_clk_i clknet_5_1__leaf_clk_i clknet_leaf_433_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_83_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10721_ _05272_ _00395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_192_4060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_4071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13440_ memory\[56\]\[28\] memory\[57\]\[28\] memory\[58\]\[28\] memory\[59\]\[28\]
+ _05711_ _03748_ _02830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09097__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10652_ memory\[51\]\[16\] _03174_ _05229_ _05236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13042__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13371_ _02762_ net58 _02382_ _02763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08844__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10583_ _05039_ memory\[50\]\[16\] _05192_ _05199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15110_ _00069_ clknet_leaf_22_clk_i memory\[42\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_88_Right_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12322_ memory\[32\]\[11\] memory\[33\]\[11\] memory\[34\]\[11\] memory\[35\]\[11\]
+ _06314_ _06454_ _06527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_1_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08452__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12228__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15041_ _00000_ clknet_leaf_438_clk_i memory\[40\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12253_ _06458_ _06459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_142_1026 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09347__I _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11204_ _05528_ _00622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12184_ _06325_ _06390_ _06391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__10954__I1 _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11135_ _03348_ memory\[58\]\[19\] _05482_ _05492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12702__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11066_ _05455_ _00557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10017_ _04884_ _00079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_97_Right_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10222__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12608__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14825_ _01864_ clknet_leaf_43_clk_i memory\[33\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_116_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_125_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08627__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12084__A2 _06283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14756_ _01795_ clknet_leaf_405_clk_i memory\[31\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11968_ _05736_ _06176_ _06177_ _06178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_15_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_173_3708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13707_ _03084_ _00771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12149__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10919_ memory\[55\]\[13\] _03165_ _05374_ _05378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14687_ _01726_ clknet_leaf_358_clk_i memory\[2\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11899_ _06109_ _06110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_129_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11053__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09088__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13638_ _05715_ _03020_ _03022_ _03024_ _03025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_89_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_27_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08835__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10892__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13569_ memory\[52\]\[30\] memory\[53\]\[30\] _05716_ _02957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11595__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_4_Left_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15308_ _00267_ clknet_leaf_258_clk_i memory\[48\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07090_ _03215_ memory\[16\]\[29\] _03251_ _03261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_2_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12139__A3 _06330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15239_ _00198_ clknet_leaf_271_clk_i memory\[46\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_131_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09800_ _04768_ _02058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13708__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12612__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07992_ _03149_ _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_5_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09193__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07706__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09012__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_163_Right_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_157_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06943_ _03162_ _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_09731_ _04731_ _02026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13195__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12847__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12698__I1 net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11228__S _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09662_ _04606_ memory\[37\]\[15\] _04689_ _04695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_2_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08613_ _04108_ _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_2_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09593_ _04658_ _01961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11027__I _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13443__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08544_ _03124_ _03225_ _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_82_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13272__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07441__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08475_ _04035_ _01466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_56_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07426_ memory\[49\]\[5\] _03319_ _03455_ _03461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10881__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11898__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08826__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07357_ _03422_ _00961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_162_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13398__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07288_ memory\[11\]\[6\] _03321_ _03379_ _03386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09027_ _04343_ _01710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10936__I1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_130_Right_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09003__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09929_ _04598_ memory\[41\]\[11\] _04836_ _04838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11138__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10042__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12940_ _05655_ _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07565__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_333_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07415__I _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output43_I net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11361__I1 _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12871_ memory\[36\]\[19\] memory\[37\]\[19\] _06447_ _02270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14610_ _01649_ clknet_leaf_81_clk_i memory\[26\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_372_clk_i clknet_5_12__leaf_clk_i clknet_leaf_372_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11822_ _06031_ _06033_ _06034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_68_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08447__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15590_ _00549_ clknet_leaf_234_clk_i memory\[57\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_29__f_clk_i clknet_2_3_0_clk_i clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12477__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09630__I _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_190_4019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14541_ _01580_ clknet_leaf_187_clk_i memory\[24\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11753_ memory\[36\]\[3\] memory\[37\]\[3\] _05733_ _05966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10704_ _05263_ _00387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13015__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_120_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14472_ _01511_ clknet_leaf_175_clk_i memory\[22\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11684_ memory\[36\]\[2\] memory\[37\]\[2\] _05733_ _05898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_387_clk_i clknet_5_6__leaf_clk_i clknet_leaf_387_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_187_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_181_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13423_ _02501_ _02813_ _02814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10635_ memory\[51\]\[8\] _03149_ _05218_ _05227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08817__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11577__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_51_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13354_ _02336_ _02738_ _02745_ _02746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_106_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08182__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10566_ _05022_ memory\[50\]\[8\] _05181_ _05190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11672__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12305_ memory\[6\]\[11\] memory\[7\]\[11\] _06431_ _06510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_106_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_310_clk_i clknet_5_11__leaf_clk_i clknet_leaf_310_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_84_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13285_ _02677_ _02678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10217__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10497_ _05153_ _00290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12236_ _06031_ _06441_ _06442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15024_ _02063_ clknet_leaf_89_clk_i memory\[3\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10927__I1 _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09793__I1 _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12167_ _06028_ _06373_ _06304_ _06374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_166_3567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11118_ _05483_ _00581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13177__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12098_ memory\[8\]\[8\] memory\[9\]\[8\] memory\[10\]\[8\] memory\[11\]\[8\] _05893_
+ _06032_ _06306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XTAP_TAPCELL_ROW_183_3892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_127_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11049_ _05026_ memory\[57\]\[10\] _05446_ _05447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput7 data_i[0] net7 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09741__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10887__S _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14808_ _01847_ clknet_leaf_68_clk_i memory\[32\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15788_ _00747_ clknet_leaf_252_clk_i net47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09540__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10686__I _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14739_ _01778_ clknet_leaf_90_clk_i memory\[30\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_143_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08260_ _03806_ memory\[17\]\[26\] _03915_ _03922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_28_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08681__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07211_ memory\[39\]\[12\] _03334_ _03330_ _03335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08191_ _03885_ _01332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12607__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07995__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07142_ _03267_ _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_15_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12860__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07073_ _03252_ _00847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12406__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_282_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09916__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09233__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08820__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13438__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11040__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09784__I1 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12342__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07795__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07975_ _03756_ memory\[12\]\[2\] _03752_ _03757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09714_ _04722_ _02018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06926_ _03149_ _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13493__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11343__I1 _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07235__I _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_87_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09645_ _04589_ memory\[37\]\[7\] _04678_ _04686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_87_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10797__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13173__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_48_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09576_ _04649_ _01953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08527_ _04063_ _01490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_65_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10854__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08458_ _03800_ memory\[20\]\[23\] _04023_ _04027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07409_ _03449_ _00986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08389_ _03990_ _01425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10420_ _05012_ memory\[48\]\[3\] _05109_ _05113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10606__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_104_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_455 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10351_ _05076_ _00221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09826__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13070_ memory\[0\]\[22\] memory\[1\]\[22\] memory\[2\]\[22\] memory\[3\]\[22\] _06709_
+ _06779_ _02466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09224__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10282_ _05030_ _00198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_148_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12021_ _06162_ _06229_ _06230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12252__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07346__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13484__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13972_ _01011_ clknet_leaf_156_clk_i memory\[49\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11334__I1 _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15711_ _00670_ clknet_leaf_334_clk_i memory\[61\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_161_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12923_ _02320_ _02321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_87_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_122_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06984__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10500__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15642_ _00601_ clknet_leaf_379_clk_i memory\[58\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08177__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12854_ _06831_ _02248_ _02250_ _02252_ _02253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_158_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11098__I0 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_85_Left_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11805_ memory\[6\]\[4\] memory\[7\]\[4\] _05706_ _06017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15573_ _00532_ clknet_leaf_160_clk_i memory\[56\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12785_ _02184_ _02185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_84_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14524_ _01563_ clknet_leaf_377_clk_i memory\[24\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11736_ _05676_ _05944_ _05946_ _05948_ _05949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08905__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07710__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14455_ _01494_ clknet_leaf_98_clk_i memory\[21\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11667_ _05651_ _05873_ _05880_ _05881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_154_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13406_ _02341_ _02796_ _05708_ _02797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10618_ _05217_ _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14386_ _01425_ clknet_leaf_139_clk_i memory\[1\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11598_ memory\[54\]\[1\] memory\[55\]\[1\] _05684_ _05813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11645__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13337_ _05777_ _02728_ _02729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10549_ _05180_ _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_109_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_168_3618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11970__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_94_Left_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09736__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13268_ _06844_ _02656_ _02658_ _02660_ _02661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_185_3932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15007_ _02046_ clknet_leaf_357_clk_i memory\[3\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11022__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_264_clk_i clknet_5_13__leaf_clk_i clknet_leaf_264_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12219_ _06149_ _06424_ _06425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13199_ memory\[4\]\[24\] memory\[5\]\[24\] _06845_ _02593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07760_ _03111_ memory\[6\]\[0\] _03639_ _03640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_279_clk_i clknet_5_12__leaf_clk_i clknet_leaf_279_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_2_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07691_ _03602_ _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_63_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11581__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09430_ _04218_ memory\[34\]\[17\] _04549_ _04557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__06894__I _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_229_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10410__S _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13227__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_202_clk_i clknet_5_30__leaf_clk_i clknet_leaf_202_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09361_ _04520_ _01867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_176_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08312_ _03949_ _01389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13721__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09292_ _04216_ memory\[32\]\[16\] _04477_ _04484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08243_ _03789_ memory\[17\]\[18\] _03904_ _03913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_8_clk_i clknet_5_5__leaf_clk_i clknet_leaf_8_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_133_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13086__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_217_clk_i clknet_5_27__leaf_clk_i clknet_leaf_217_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08174_ _03876_ _01324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08614__I _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07125_ _03281_ _00870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_166_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11261__I0 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11961__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07056_ _03243_ _00839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08550__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13168__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07768__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07958_ _03218_ memory\[19\]\[30\] _03710_ _03744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09381__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06909_ net33 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07889_ _03707_ _01208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_104_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09628_ _04676_ _01978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07940__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09559_ _04639_ memory\[35\]\[31\] _04574_ _04640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_100_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_65_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10827__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_80_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12570_ memory\[48\]\[15\] memory\[49\]\[15\] memory\[50\]\[15\] memory\[51\]\[15\]
+ _06699_ _06150_ _06771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08725__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09693__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12755__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11521_ _05683_ _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_80_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11452_ _05667_ _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14240_ _01279_ clknet_leaf_278_clk_i memory\[15\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09445__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10403_ _05103_ _00246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14171_ _01210_ clknet_leaf_393_clk_i memory\[7\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11383_ _03323_ memory\[62\]\[7\] _05616_ _05624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12744__A3 _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09556__S _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13122_ _02516_ _02517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10334_ _05065_ _00215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08460__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11004__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13053_ memory\[62\]\[22\] memory\[63\]\[22\] _02448_ _02449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_178_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06979__I net20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10265_ _05018_ memory\[46\]\[6\] _05006_ _05019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07076__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12004_ _05660_ _06212_ _06001_ _06213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10196_ _04593_ memory\[45\]\[9\] _04969_ _04979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_180_3840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13457__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11307__I1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07804__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13955_ _00994_ clknet_leaf_334_clk_i memory\[49\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08184__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11326__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_230_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12906_ _02303_ _02304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__10230__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13209__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13886_ _00925_ clknet_leaf_309_clk_i memory\[11\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07931__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_57_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15625_ _00584_ clknet_leaf_233_clk_i memory\[58\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12837_ _06467_ _02228_ _02236_ _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_68_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15556_ _00515_ clknet_leaf_319_clk_i memory\[56\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12768_ memory\[62\]\[18\] memory\[63\]\[18\] _06557_ _02168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_56_344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14507_ _01546_ clknet_leaf_197_clk_i memory\[23\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11719_ _05767_ _05925_ _05932_ _05933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__12157__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12983__A3 _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15487_ _00446_ clknet_leaf_331_clk_i memory\[54\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11061__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12699_ _02100_ _00747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14438_ _01477_ clknet_leaf_188_clk_i memory\[21\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput10 data_i[12] net10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput21 data_i[22] net21 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xinput32 data_i[3] net32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14369_ _01408_ clknet_leaf_340_clk_i memory\[1\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11943__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_23_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08930_ _04292_ _01664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06889__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13240__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08861_ _04193_ memory\[26\]\[5\] _04250_ _04256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_36_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07812_ _03203_ memory\[6\]\[25\] _03661_ _03667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08792_ _04210_ memory\[25\]\[13\] _04204_ _04211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13448__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07743_ _03630_ _01139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08175__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12120__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07674_ _03200_ memory\[10\]\[24\] _03589_ _03594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_141_clk_i clknet_5_19__leaf_clk_i clknet_leaf_141_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_95_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_95_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_176_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09413_ _04201_ memory\[34\]\[9\] _04538_ _04548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13451__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10809__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09344_ _04511_ _01859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13620__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09675__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09275_ _04199_ memory\[32\]\[8\] _04466_ _04475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_156_clk_i clknet_5_24__leaf_clk_i clknet_leaf_156_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_63_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_432_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08226_ _03892_ _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_28_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12806__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11234__I0 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08157_ _03867_ _01316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07108_ _03272_ _00862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08088_ _03818_ _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08280__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08650__I1 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07039_ _03234_ _00831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10315__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10050_ _04583_ memory\[43\]\[4\] _04897_ _04902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_73_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13439__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07624__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11146__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_109_clk_i clknet_5_22__leaf_clk_i clknet_leaf_109_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13740_ _03359_ memory\[9\]\[24\] _03097_ _03102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10050__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08519__I _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10952_ memory\[55\]\[29\] _03214_ _05385_ _05395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_27_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13671_ _03057_ _03058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_97_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10985__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10883_ _05066_ memory\[54\]\[29\] _05348_ _05358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_94_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15410_ _00369_ clknet_leaf_153_clk_i memory\[51\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12622_ _06822_ _00746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09666__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_159_Left_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_66_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15341_ _00300_ clknet_leaf_251_clk_i memory\[4\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12553_ _06484_ _06754_ _06755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_156_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_156_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11504_ _05683_ _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_81_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15272_ _00231_ clknet_leaf_272_clk_i memory\[47\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09418__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12484_ _06686_ _00744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12178__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14223_ _01262_ clknet_leaf_197_clk_i memory\[12\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11435_ _03450_ _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_134_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13470__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09286__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14154_ _01193_ clknet_leaf_221_clk_i memory\[7\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08190__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11366_ _05614_ _00698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11829__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_120_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13105_ _05667_ _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_10317_ _03196_ _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_120_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_130_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14085_ _01124_ clknet_leaf_303_clk_i memory\[63\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11297_ _05577_ _00666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_168_Left_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13036_ memory\[24\]\[21\] memory\[25\]\[21\] memory\[26\]\[21\] memory\[27\]\[21\]
+ _02363_ _06611_ _02433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_10248_ _05007_ _00187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13536__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10179_ _04970_ _00155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07534__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13525__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10959__I _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14987_ _02026_ clknet_leaf_43_clk_i memory\[38\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_381_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13938_ _00977_ clknet_leaf_123_clk_i memory\[8\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07904__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13869_ _00908_ clknet_leaf_263_clk_i memory\[39\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_177_Left_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13271__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_73_clk_i clknet_5_16__leaf_clk_i clknet_leaf_73_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15608_ _00567_ clknet_leaf_269_clk_i memory\[57\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07390_ _03194_ memory\[8\]\[22\] _03437_ _03440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08365__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13602__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15539_ _00498_ clknet_leaf_153_clk_i memory\[55\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_09060_ _04361_ _01725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09409__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_88_clk_i clknet_5_20__leaf_clk_i clknet_leaf_88_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12169__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08011_ _03168_ _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_128_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11216__I0 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11916__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_186_Left_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_38_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_11_clk_i clknet_5_5__leaf_clk_i clknet_leaf_11_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_38_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10135__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09962_ _04631_ memory\[41\]\[27\] _04847_ _04855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13669__A1 _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09924__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08913_ _04245_ memory\[26\]\[30\] _04249_ _04283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_55_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09893_ _04818_ _00021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08396__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08844_ _04245_ memory\[25\]\[30\] _04182_ _04246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_26_clk_i clknet_5_4__leaf_clk_i clknet_leaf_26_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08775_ _03149_ _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_169_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08148__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07726_ _03621_ _01131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09896__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_126_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07657_ _03175_ memory\[10\]\[16\] _03578_ _03585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11998__A4 _06207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_0_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07588_ _03175_ memory\[0\]\[16\] _03541_ _03548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09327_ _04181_ memory\[33\]\[0\] _04502_ _04503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08320__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_11_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10958__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09258_ _04465_ _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_185_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08209_ _03895_ _01340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10109__I _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09189_ _03306_ _03855_ _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_161_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_177_Right_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_151_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11220_ _03365_ memory\[5\]\[27\] _05529_ _05537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07619__S _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08623__I1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12580__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_112_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11151_ _05500_ _00597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10102_ _04635_ memory\[43\]\[29\] _04919_ _04929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11082_ _05060_ memory\[57\]\[26\] _05457_ _05464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12332__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14910_ _01949_ clknet_leaf_436_clk_i memory\[36\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10033_ _04892_ _00087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10194__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07354__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14841_ _01880_ clknet_leaf_70_clk_i memory\[33\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14772_ _01811_ clknet_leaf_90_clk_i memory\[31\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11984_ memory\[30\]\[6\] memory\[31\]\[6\] _06193_ _06194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12191__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13723_ _03342_ memory\[9\]\[16\] _03086_ _03093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10935_ _05386_ _00495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11604__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06992__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09639__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13654_ _03114_ _03033_ _03040_ _03041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_112_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_175_3750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10866_ _05349_ _00463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_184_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12605_ memory\[28\]\[15\] memory\[29\]\[15\] _06604_ _06806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_54_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13104__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13585_ _02972_ _02973_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_112_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08311__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10797_ _05047_ memory\[53\]\[20\] _05312_ _05313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15324_ _00283_ clknet_leaf_368_clk_i memory\[4\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_171_3658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_42_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12536_ memory\[40\]\[14\] memory\[41\]\[14\] memory\[42\]\[14\] memory\[43\]\[14\]
+ _06186_ _06326_ _06738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_87_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_171_3669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08913__S _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_152_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_132_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_328_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15255_ _00214_ clknet_leaf_41_clk_i memory\[46\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12467_ memory\[28\]\[13\] memory\[29\]\[13\] _06604_ _06670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_144_Right_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14206_ _01245_ clknet_leaf_373_clk_i memory\[12\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11418_ _05642_ _00722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15186_ _00145_ clknet_leaf_14_clk_i memory\[44\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12398_ _06445_ _06593_ _06601_ _06602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__12571__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14137_ _01176_ clknet_leaf_142_clk_i memory\[6\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11349_ memory\[61\]\[23\] _03196_ _05602_ _05606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14068_ _01107_ clknet_leaf_129_clk_i memory\[10\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11757__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13019_ memory\[38\]\[21\] memory\[39\]\[21\] _06728_ _02416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06890_ net39 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_146_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09543__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08560_ _03766_ memory\[22\]\[7\] _04073_ _04081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07511_ memory\[59\]\[12\] _03334_ _03504_ _03507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08491_ _04044_ _01473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_18_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07998__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08550__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07442_ _03469_ _00999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08095__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07373_ _03169_ memory\[8\]\[14\] _03426_ _03431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09112_ _04388_ _01750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08823__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_96_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09043_ _04239_ memory\[28\]\[27\] _04344_ _04352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07439__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_111_Right_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_92_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12562__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09654__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07238__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09945_ _04614_ memory\[41\]\[19\] _04836_ _04846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08369__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11983__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_70_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09876_ _04809_ _00013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07174__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08827_ _04234_ _01619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08758_ _04187_ memory\[25\]\[2\] _04183_ _04188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09869__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07902__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07709_ _03612_ _01123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_277_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08689_ _03758_ memory\[24\]\[3\] _04146_ _04150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10720_ _05039_ memory\[52\]\[16\] _05265_ _05272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_192_4061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_4072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_136_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10651_ _05235_ _00362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13370_ _02716_ _02731_ _02746_ _02761_ _02762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_24_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10100__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10582_ _05198_ _00330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08733__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12321_ _06450_ _06525_ _06177_ _06526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_133_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12228__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15040_ _02079_ clknet_leaf_438_clk_i memory\[40\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_106_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12252_ memory\[44\]\[10\] memory\[45\]\[10\] _06319_ _06458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11203_ _03348_ memory\[5\]\[19\] _05518_ _05528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11987__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12183_ memory\[40\]\[9\] memory\[41\]\[9\] memory\[42\]\[9\] memory\[43\]\[9\] _06186_
+ _06326_ _06390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_102_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11134_ _05491_ _00589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11065_ _05043_ memory\[57\]\[18\] _05446_ _05455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10503__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06987__I net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07084__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07032__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10016_ _04616_ memory\[42\]\[20\] _04883_ _04884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14824_ _01863_ clknet_leaf_45_clk_i memory\[33\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07812__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_98_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14755_ _01794_ clknet_leaf_410_clk_i memory\[31\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11967_ _05686_ _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08532__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11334__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13706_ _03325_ memory\[9\]\[8\] _03075_ _03084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10918_ _05377_ _00487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14686_ _01725_ clknet_leaf_359_clk_i memory\[2\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_156_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11898_ memory\[44\]\[5\] memory\[45\]\[5\] _05749_ _06109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11419__I0 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13637_ _05724_ _03023_ _03024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10849_ _05340_ _00455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13568_ _05700_ _02951_ _02953_ _02955_ _02956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_70_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_14_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15307_ _00266_ clknet_leaf_234_clk_i memory\[48\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12519_ _03747_ _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10642__I1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13499_ memory\[60\]\[29\] memory\[61\]\[29\] _05702_ _02888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15238_ _00197_ clknet_leaf_271_clk_i memory\[46\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12139__A4 _06346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_188_3985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15169_ _00128_ clknet_leaf_421_clk_i memory\[44\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_188_3996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07991_ _03767_ _01250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09730_ _04606_ memory\[38\]\[15\] _04725_ _04731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10158__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06942_ net10 _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_158_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09661_ _04694_ _01993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_105_Left_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_2_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08612_ _03225_ _03306_ _04108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_09592_ _04604_ memory\[36\]\[14\] _04653_ _04658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08543_ _04071_ _01498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07326__I1 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11244__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11902__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08474_ _03816_ memory\[20\]\[31\] _04000_ _04035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10330__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07425_ _03460_ _00991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09649__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07356_ _03144_ memory\[8\]\[6\] _03415_ _03422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12783__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10633__I1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07287_ _03385_ _00928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13407__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09026_ _04222_ memory\[28\]\[19\] _04333_ _04343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_851 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12535__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11969__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12803__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11927__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_141_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11419__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09928_ _04837_ _00037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10149__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09859_ _04595_ memory\[40\]\[10\] _04800_ _04801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_99_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13634__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_107_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12870_ _06428_ _02261_ _02268_ _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_107_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12146__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07632__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11821_ memory\[8\]\[4\] memory\[9\]\[4\] memory\[10\]\[4\] memory\[11\]\[4\] _05893_
+ _06032_ _06033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_139_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11154__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14540_ _01579_ clknet_leaf_188_clk_i memory\[24\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11752_ _05699_ _05957_ _05964_ _05965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_166_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10321__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10703_ _05022_ memory\[52\]\[8\] _05254_ _05263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14471_ _01510_ clknet_leaf_171_clk_i memory\[22\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_120_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10993__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11683_ _05699_ _05888_ _05896_ _05897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_138_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13422_ memory\[24\]\[27\] memory\[25\]\[27\] memory\[26\]\[27\] memory\[27\]\[27\]
+ _02363_ _02502_ _02813_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__09559__S _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10634_ _05226_ _00354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12774__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13353_ _02209_ _02740_ _02742_ _02744_ _02745_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10565_ _05189_ _00322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12304_ _06508_ _06509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_20_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13284_ memory\[44\]\[25\] memory\[45\]\[25\] _02210_ _02677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10496_ _05020_ memory\[4\]\[7\] _05145_ _05153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_51_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15023_ _02062_ clknet_leaf_168_clk_i memory\[3\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12235_ memory\[8\]\[10\] memory\[9\]\[10\] memory\[10\]\[10\] memory\[11\]\[10\]
+ _05893_ _06032_ _06441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__10388__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09294__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12166_ memory\[14\]\[9\] memory\[15\]\[9\] _06302_ _06373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_166_3568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_166_3579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12512__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11117_ _03329_ memory\[58\]\[10\] _05482_ _05483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12097_ _06028_ _06303_ _06304_ _06305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_183_3893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07005__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_127_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11048_ _05434_ _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
Xinput8 data_i[10] net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__13544__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10560__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07542__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14807_ _01846_ clknet_leaf_73_clk_i memory\[32\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15787_ _00746_ clknet_leaf_254_clk_i net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08505__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12999_ _06838_ _02395_ _02396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_8_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14738_ _01777_ clknet_leaf_88_clk_i memory\[30\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10312__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_131_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14669_ _01708_ clknet_leaf_184_clk_i memory\[28\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07210_ _03162_ _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08190_ _03804_ memory\[29\]\[25\] _03879_ _03885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08373__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11798__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07141_ _03289_ _00878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10408__S _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12860__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_41_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07072_ _03187_ memory\[16\]\[20\] _03251_ _03252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_225_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12517__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13719__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12623__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10379__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07717__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13190__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_432_clk_i clknet_5_1__leaf_clk_i clknet_leaf_432_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10143__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07974_ _03131_ _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_113_Left_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09713_ _04589_ memory\[38\]\[7\] _04714_ _04722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06925_ net37 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09697__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09644_ _04685_ _01985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_87_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08548__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09575_ _04587_ memory\[36\]\[6\] _04642_ _04649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08526_ _03800_ memory\[21\]\[23\] _04059_ _04063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08457_ _04026_ _01457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_122_Left_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_136_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11702__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09379__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07408_ _03221_ memory\[8\]\[31\] _03414_ _03449_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08388_ _03798_ memory\[1\]\[22\] _03987_ _03990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13202__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11803__I0 memory\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07339_ _03412_ _00953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10318__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10350_ _05010_ memory\[47\]\[2\] _05073_ _05076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09009_ _04334_ _01701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10281_ _05029_ memory\[46\]\[11\] _05027_ _05030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13181__A1 _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12020_ memory\[0\]\[7\] memory\[1\]\[7\] memory\[2\]\[7\] memory\[3\]\[7\] _06020_
+ _06090_ _06229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_108_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_148_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_131_Left_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08983__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10790__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09842__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_427_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13971_ _01010_ clknet_leaf_157_clk_i memory\[49\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08735__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07538__I1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13364__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15710_ _00669_ clknet_leaf_334_clk_i memory\[61\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_161_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12922_ memory\[4\]\[20\] memory\[5\]\[20\] _06845_ _02320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08458__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10542__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07362__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12119__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15641_ _00600_ clknet_leaf_268_clk_i memory\[58\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12853_ _06838_ _02251_ _02252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_122_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11804_ _06015_ _06016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15572_ _00531_ clknet_leaf_166_clk_i memory\[56\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12784_ memory\[4\]\[18\] memory\[5\]\[18\] _06845_ _02184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_174_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_140_Left_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09160__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14523_ _01562_ clknet_leaf_398_clk_i memory\[23\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11735_ _05690_ _05947_ _05948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14454_ _01493_ clknet_leaf_93_clk_i memory\[21\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_148_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11666_ _05676_ _05875_ _05877_ _05879_ _05880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_154_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13405_ memory\[38\]\[27\] memory\[39\]\[27\] _05662_ _02796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10617_ _05216_ _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_14385_ _01424_ clknet_leaf_109_clk_i memory\[1\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12507__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10228__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11597_ _05811_ _05812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_141_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13336_ memory\[8\]\[26\] memory\[9\]\[26\] memory\[10\]\[26\] memory\[11\]\[26\]
+ _02473_ _05779_ _02728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_51_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08921__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10548_ _03451_ _03565_ _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_168_3608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_168_3619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13267_ _06851_ _02659_ _02660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_62_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10479_ _05143_ _00282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13172__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15006_ _02045_ clknet_leaf_357_clk_i memory\[3\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07226__I0 memory\[39\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12218_ memory\[48\]\[10\] memory\[49\]\[10\] memory\[50\]\[10\] memory\[51\]\[10\]
+ _06010_ _06150_ _06424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_13198_ _02302_ _02584_ _02591_ _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_20_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11059__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_99_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12149_ memory\[52\]\[9\] memory\[53\]\[9\] _06143_ _06356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10898__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07690_ _03306_ _03490_ _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_154_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11581__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09360_ _04216_ memory\[33\]\[16\] _04513_ _04520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07071__I _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_19_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08311_ _03789_ memory\[18\]\[18\] _03940_ _03949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_192_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09291_ _04483_ _01834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11522__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_43_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09199__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08242_ _03912_ _01356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_62_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13086__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08173_ _03787_ memory\[29\]\[17\] _03868_ _03876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12202__A3 _06393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11321__I _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07124_ _03160_ memory\[13\]\[11\] _03279_ _03281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09927__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_376_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07055_ _03163_ memory\[16\]\[12\] _03240_ _03243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11961__A2 _06170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_371_clk_i clknet_5_9__leaf_clk_i clknet_leaf_371_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13163__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07217__I0 memory\[39\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08965__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12910__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12761__I1 net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_89_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09662__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input35_I data_i[6] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07957_ _03743_ _01240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_386_clk_i clknet_5_6__leaf_clk_i clknet_leaf_386_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_143_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13184__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06908_ _03136_ _00798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08278__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10524__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07888_ _03215_ memory\[7\]\[29\] _03697_ _03707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09461__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09627_ _04639_ memory\[36\]\[31\] _04641_ _04676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09558_ _03220_ _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_100_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07910__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08509_ _03783_ memory\[21\]\[15\] _04048_ _04054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09489_ _04592_ _01923_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_80_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11520_ _05659_ _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_65_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_324_clk_i clknet_5_10__leaf_clk_i clknet_leaf_324_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_0_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12729__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_4011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11451_ _03117_ _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10048__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11231__I _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10402_ _05062_ memory\[47\]\[27\] _05095_ _05103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14170_ _01209_ clknet_leaf_393_clk_i memory\[7\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08741__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11382_ _05623_ _00705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13121_ memory\[60\]\[23\] memory\[61\]\[23\] _02164_ _02516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_339_clk_i clknet_5_9__leaf_clk_i clknet_leaf_339_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_46_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10333_ _05064_ memory\[46\]\[28\] _05048_ _05065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_115_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07208__I0 memory\[39\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13052_ _05661_ _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_10264_ _03143_ _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_44_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08956__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12003_ memory\[62\]\[7\] memory\[63\]\[7\] _05868_ _06212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_163_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10195_ _04978_ _00163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10763__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08708__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13954_ _00993_ clknet_leaf_315_clk_i memory\[49\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10511__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06995__I net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_22__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08188__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10515__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07092__S _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09381__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12905_ memory\[60\]\[20\] memory\[61\]\[20\] _02164_ _02303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13885_ _00924_ clknet_leaf_288_clk_i memory\[11\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12011__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12836_ _06476_ _02230_ _02232_ _02235_ _02236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_124_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15624_ _00583_ clknet_leaf_234_clk_i memory\[58\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07820__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09133__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_13__f_clk_i clknet_2_1_0_clk_i clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_189_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12968__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15555_ _00514_ clknet_leaf_321_clk_i memory\[56\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12767_ _05659_ _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14506_ _01545_ clknet_leaf_173_clk_i memory\[23\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11718_ _05783_ _05927_ _05929_ _05931_ _05932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__11640__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15486_ _00445_ clknet_leaf_331_clk_i memory\[54\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12698_ _02099_ net47 _06491_ _02100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14437_ _01476_ clknet_leaf_375_clk_i memory\[21\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11649_ _05818_ _05833_ _05848_ _05863_ _05864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
Xinput11 data_i[13] net11 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput22 data_i[23] net22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__13393__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput33 data_i[4] net33 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09747__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14368_ _01407_ clknet_leaf_341_clk_i memory\[1\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13269__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13319_ memory\[54\]\[26\] memory\[55\]\[26\] _02312_ _02711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10980__I _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14299_ _01338_ clknet_leaf_1_clk_i memory\[29\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09546__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12579__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13240__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08860_ _04255_ _01631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09482__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07811_ _03666_ _01171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_36_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08791_ _03165_ _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_58_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07742_ _03200_ memory\[63\]\[24\] _03625_ _03630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12120__A2 _06327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07673_ _03593_ _01106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_149_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13732__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09412_ _04547_ _01891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06886__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08826__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12959__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09343_ _04199_ memory\[33\]\[8\] _04502_ _04511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_158_Right_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07686__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09274_ _04474_ _01826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11631__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08225_ _03903_ _01348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12806__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08156_ _03770_ memory\[29\]\[9\] _03857_ _03867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07107_ _03135_ memory\[13\]\[3\] _03268_ _03272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10890__I _05361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08087_ _03829_ _01284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10993__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07177__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_122_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07038_ _03138_ memory\[16\]\[4\] _03229_ _03234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_77_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11698__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12811__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10745__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08989_ _04185_ memory\[28\]\[1\] _04322_ _04324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13439__A2 _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11427__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10951_ _05394_ _00503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11170__I0 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13642__S _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10130__I _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11870__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13670_ memory\[28\]\[31\] memory\[29\]\[31\] _02495_ _03057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10882_ _05357_ _00471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09115__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07640__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12621_ _06821_ net46 _06491_ _06822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_263_clk_i clknet_5_13__leaf_clk_i clknet_leaf_263_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_47_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_125_Right_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_108_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15340_ _00299_ clknet_leaf_252_clk_i memory\[4\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12552_ memory\[16\]\[14\] memory\[17\]\[14\] memory\[18\]\[14\] memory\[19\]\[14\]
+ _06342_ _06485_ _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__11622__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11503_ _05681_ _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_136_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15271_ _00230_ clknet_leaf_271_clk_i memory\[47\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12483_ _06685_ net44 _06491_ _06686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_117_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14222_ _01261_ clknet_leaf_195_clk_i memory\[12\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09567__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11434_ _05650_ _00730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_278_clk_i clknet_5_12__leaf_clk_i clknet_leaf_278_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_151_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13089__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13470__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14153_ _01192_ clknet_leaf_221_clk_i memory\[7\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11365_ memory\[61\]\[31\] _03220_ _05579_ _05614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_162_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13127__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13104_ _02498_ _02499_ _02086_ _02500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10316_ _05053_ _00209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14084_ _01123_ clknet_leaf_305_clk_i memory\[63\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11296_ _03373_ memory\[60\]\[31\] _05542_ _05577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_201_clk_i clknet_5_30__leaf_clk_i clknet_leaf_201_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_123_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08929__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13035_ _06607_ _02431_ _02086_ _02432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__11689__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10247_ _05004_ memory\[46\]\[0\] _05006_ _05007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07601__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10178_ _04573_ memory\[45\]\[0\] _04969_ _04970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_7_clk_i clknet_5_5__leaf_clk_i clknet_leaf_7_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_156_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_216_clk_i clknet_5_27__leaf_clk_i clknet_leaf_216_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14986_ _02025_ clknet_leaf_43_clk_i memory\[38\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_324_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09354__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13937_ _00976_ clknet_leaf_123_clk_i memory\[8\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_187_954 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13868_ _00907_ clknet_leaf_258_clk_i memory\[39\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07550__S _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12819_ _02216_ _02218_ _02219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15607_ _00566_ clknet_leaf_159_clk_i memory\[57\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13799_ _00838_ clknet_leaf_204_clk_i memory\[16\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11072__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07668__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15538_ _00497_ clknet_leaf_153_clk_i memory\[55\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15469_ _00428_ clknet_leaf_289_clk_i memory\[53\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08010_ _03780_ _01256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12169__A2 _06375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08381__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_142_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08093__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10416__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13118__A1 _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_38_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09961_ _04854_ _00053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07840__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13727__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08912_ _04282_ _01656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09892_ _04629_ memory\[40\]\[26\] _04811_ _04818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07725__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08843_ _03217_ _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_85_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08774_ _04198_ _01602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_26_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09345__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07725_ _03175_ memory\[63\]\[16\] _03614_ _03621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11152__I0 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07656_ _03584_ _01098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11852__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08556__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07460__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_0_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12078__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07587_ _03547_ _01066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07659__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09326_ _04501_ _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_35_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_11_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_63_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09257_ net73 _03305_ _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_8_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_173_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08208_ _03754_ memory\[17\]\[1\] _03893_ _03895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09387__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09188_ _04428_ _01786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_151_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08139_ _03858_ _01307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08084__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10966__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13109__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09820__I1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_75_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_273_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11150_ _03363_ memory\[58\]\[26\] _05493_ _05500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_112_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10101_ _04928_ _00119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11081_ _05463_ _00564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10718__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output66_I net66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09584__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10032_ _04633_ memory\[42\]\[28\] _04883_ _04892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14840_ _01879_ clknet_leaf_69_clk_i memory\[33\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09850__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14771_ _01810_ clknet_leaf_90_clk_i memory\[31\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11983_ _05683_ _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13722_ _03092_ _00778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_98_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07898__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12191__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10934_ memory\[55\]\[20\] _03186_ _05385_ _05386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08466__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_158_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12496__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_112_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13653_ _05768_ _03035_ _03037_ _03039_ _03040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_156_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10865_ _05047_ memory\[54\]\[20\] _05348_ _05349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_175_3740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_27_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13140__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12604_ _06445_ _06797_ _06804_ _06805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_183_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13584_ memory\[12\]\[30\] memory\[13\]\[30\] _05769_ _02972_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10796_ _05289_ _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_82_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15323_ _00282_ clknet_leaf_374_clk_i memory\[48\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12535_ _06322_ _06736_ _06461_ _06737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_171_3659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15254_ _00213_ clknet_leaf_41_clk_i memory\[46\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12466_ _06445_ _06661_ _06668_ _06669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_151_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07027__A1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14205_ _01244_ clknet_leaf_270_clk_i memory\[12\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11417_ _03357_ memory\[62\]\[23\] _05638_ _05642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12515__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10236__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15185_ _00144_ clknet_leaf_14_clk_i memory\[44\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_2_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12397_ _06318_ _06595_ _06598_ _06600_ _06601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
Xclkbuf_leaf_140_clk_i clknet_5_22__leaf_clk_i clknet_leaf_140_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09096__I _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14136_ _01175_ clknet_leaf_142_clk_i memory\[6\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11348_ _05605_ _00689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07822__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14067_ _01106_ clknet_leaf_120_clk_i memory\[10\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11279_ _05568_ _00657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13520__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09575__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13018_ _02414_ _02415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__13371__I1 net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11757__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_155_clk_i clknet_5_24__leaf_clk_i clknet_leaf_155_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11067__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09327__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14969_ _02008_ clknet_leaf_14_clk_i memory\[37\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07510_ _03506_ _01030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08490_ _03764_ memory\[21\]\[6\] _04037_ _04044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07280__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07441_ memory\[49\]\[12\] _03334_ _03466_ _03469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13587__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07372_ _03430_ _00968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_169_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09111_ _04239_ memory\[2\]\[27\] _04380_ _04388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13339__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09042_ _04351_ _01717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_53_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1053 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12011__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13030__B _02424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_108_clk_i clknet_5_20__leaf_clk_i clknet_leaf_108_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09935__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09944_ _04845_ _00045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12361__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13511__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09875_ _04612_ memory\[40\]\[18\] _04800_ _04809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11373__I0 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08826_ _04233_ memory\[25\]\[24\] _04225_ _04234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09670__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08757_ _03131_ _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11125__I0 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11705__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07708_ _03150_ memory\[63\]\[8\] _03603_ _03612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08286__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08688_ _04149_ _01565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_184_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07639_ _03575_ _01090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11504__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10650_ memory\[51\]\[15\] _03171_ _05229_ _05235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09309_ _04233_ memory\[32\]\[24\] _04488_ _04493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_153_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10581_ _05037_ memory\[50\]\[15\] _05192_ _05198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12320_ memory\[38\]\[11\] memory\[39\]\[11\] _06039_ _06525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08813__I _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12251_ _06446_ _06449_ _06452_ _06456_ _06457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10056__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11202_ _05527_ _00621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07804__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12553__A2 _06754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11987__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12182_ _06322_ _06388_ _05757_ _06389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_11133_ _03346_ memory\[58\]\[18\] _05482_ _05491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07280__I1 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_72_clk_i clknet_5_16__leaf_clk_i clknet_leaf_72_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07365__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13502__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11064_ _05454_ _00556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10015_ _04860_ _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_129_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09309__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_87_clk_i clknet_5_20__leaf_clk_i clknet_leaf_87_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_192_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14823_ _01862_ clknet_leaf_50_clk_i memory\[33\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08196__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11966_ memory\[38\]\[6\] memory\[39\]\[6\] _06039_ _06176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14754_ _01793_ clknet_leaf_410_clk_i memory\[31\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13705_ _03083_ _00770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10917_ memory\[55\]\[12\] _03162_ _05374_ _05377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_15_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14685_ _01724_ clknet_leaf_377_clk_i memory\[2\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_10_clk_i clknet_5_5__leaf_clk_i clknet_leaf_10_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_17_Left_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11897_ _05732_ _06103_ _06105_ _06107_ _06108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_50_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13636_ memory\[48\]\[31\] memory\[49\]\[31\] memory\[50\]\[31\] memory\[51\]\[31\]
+ _05725_ _05726_ _03023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_132_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10848_ _05031_ memory\[54\]\[12\] _05337_ _05340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12446__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13567_ _05710_ _02954_ _02955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10779_ _05303_ _00422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12518_ _05689_ _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_25_clk_i clknet_5_4__leaf_clk_i clknet_leaf_25_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_82_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15306_ _00265_ clknet_leaf_235_clk_i memory\[48\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_48_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13498_ _02887_ _00759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_42_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12449_ _06031_ _06651_ _06652_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15237_ _00196_ clknet_leaf_404_clk_i memory\[46\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_26_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_125_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09755__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15168_ _00127_ clknet_leaf_422_clk_i memory\[44\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_188_3986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_26_Left_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_188_3997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13277__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14119_ _01158_ clknet_leaf_222_clk_i memory\[6\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12181__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_169_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15099_ _00058_ clknet_leaf_443_clk_i memory\[41\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07990_ _03766_ memory\[12\]\[7\] _03752_ _03767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12927__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06941_ _03161_ _00806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_157_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08220__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09660_ _04604_ memory\[37\]\[14\] _04689_ _04694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08611_ _04107_ _01530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09591_ _04657_ _01960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_221_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08542_ _03816_ memory\[21\]\[31\] _04036_ _04071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11807__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09720__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11902__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08473_ _04034_ _01465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13740__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07424_ memory\[49\]\[4\] _03317_ _03455_ _03460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07355_ _03421_ _00960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_162_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10094__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07286_ memory\[11\]\[5\] _03319_ _03379_ _03385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13407__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09025_ _04342_ _01709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12535__A2 _06736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11969__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07411__A1 _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10604__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09927_ _04595_ memory\[41\]\[10\] _04836_ _04837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12838__A3 _02221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09858_ _04788_ _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_77_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_146_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08809_ _03183_ _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_107_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09789_ memory\[3\]\[10\] _03155_ _04762_ _04763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11820_ _03747_ _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12146__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07712__I _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09711__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11751_ _05715_ _05959_ _05961_ _05963_ _05964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_178_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10702_ _05262_ _00386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14470_ _01509_ clknet_leaf_172_clk_i memory\[22\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_139_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11682_ _05715_ _05890_ _05892_ _05895_ _05896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_181_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13421_ _02498_ _02811_ _05665_ _02812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08278__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10633_ memory\[51\]\[7\] _03146_ _05218_ _05226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11026__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11657__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11170__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_423_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13352_ _02216_ _02743_ _02744_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10564_ _05020_ memory\[50\]\[7\] _05181_ _05189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12303_ memory\[4\]\[11\] memory\[5\]\[11\] _06156_ _06508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_162_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12065__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13283_ _02337_ _02671_ _02673_ _02675_ _02676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_20_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10495_ _05152_ _00289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15022_ _02061_ clknet_leaf_169_clk_i memory\[3\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09575__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12234_ _06028_ _06439_ _06304_ _06440_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_32_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_170_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12165_ _06371_ _06372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_20_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_166_3569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_9_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12909__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11116_ _05470_ _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_12096_ _05664_ _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_183_3894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11047_ _05445_ _00548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08202__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08919__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__09950__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput9 data_i[11] net9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_56_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11345__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14806_ _01845_ clknet_leaf_70_clk_i memory\[32\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15786_ _00745_ clknet_leaf_254_clk_i net45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1063 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12998_ memory\[48\]\[21\] memory\[49\]\[21\] memory\[50\]\[21\] memory\[51\]\[21\]
+ _06699_ _06839_ _02395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_19_1160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14737_ _01776_ clknet_leaf_90_clk_i memory\[30\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_52_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12462__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11949_ _05659_ _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13560__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_89_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14668_ _01707_ clknet_leaf_183_clk_i memory\[28\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_95_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13619_ _05760_ _03006_ _03007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_171_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14599_ _01638_ clknet_leaf_179_clk_i memory\[26\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11080__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09549__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07140_ _03184_ memory\[13\]\[19\] _03279_ _03289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_41_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07071_ _03228_ _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07492__I1 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09485__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12073__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08441__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10424__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07973_ _03755_ _01244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09712_ _04721_ _02017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06924_ _03148_ _00802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13573__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08829__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09697__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12859__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11763__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09643_ _04587_ memory\[37\]\[6\] _04678_ _04685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09941__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11255__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_372_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09574_ _04648_ _01952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08525_ _04062_ _01489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11887__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_65_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08456_ _03798_ memory\[20\]\[22\] _04023_ _04026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08564__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_82_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07407_ _03448_ _00985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08387_ _03989_ _01424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10067__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07338_ memory\[11\]\[30\] _03371_ _03378_ _03412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_122_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07269_ memory\[39\]\[31\] _03373_ _03308_ _03374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12814__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09008_ _04203_ memory\[28\]\[10\] _04333_ _04334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09395__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07908__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11938__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10280_ _03159_ _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_44_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13181__A2 _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13308__I1 net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08739__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13970_ _01009_ clknet_leaf_161_clk_i memory\[49\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12769__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_12__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12921_ _03114_ _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12692__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12119__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15640_ _00599_ clknet_leaf_266_clk_i memory\[58\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12852_ memory\[48\]\[19\] memory\[49\]\[19\] memory\[50\]\[19\] memory\[51\]\[19\]
+ _06699_ _06839_ _02251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_122_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11803_ memory\[4\]\[4\] memory\[5\]\[4\] _05702_ _06015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08499__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15571_ _00530_ clknet_leaf_165_clk_i memory\[56\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12783_ _06411_ _02174_ _02182_ _02183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA_clkbuf_leaf_117_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_56_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13380__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11734_ memory\[48\]\[3\] memory\[49\]\[3\] memory\[50\]\[3\] memory\[51\]\[3\] _05692_
+ _05694_ _05947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_14522_ _01561_ clknet_leaf_398_clk_i memory\[23\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_166_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08474__S _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_3_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14453_ _01492_ clknet_leaf_100_clk_i memory\[21\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11665_ _05690_ _05878_ _05879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10509__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10058__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09999__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10616_ _03376_ _03451_ _05216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_13404_ _02794_ _02795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_14384_ _01423_ clknet_leaf_109_clk_i memory\[1\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_919 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08273__I _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11596_ memory\[52\]\[1\] memory\[53\]\[1\] _05678_ _05811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13335_ _05772_ _02726_ _02195_ _02727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_40_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10547_ _05179_ _00314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10308__I _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07474__I1 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12724__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_168_3609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07818__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13266_ memory\[0\]\[25\] memory\[1\]\[25\] memory\[2\]\[25\] memory\[3\]\[25\] _05784_
+ _03226_ _02659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10478_ _05070_ memory\[48\]\[31\] _05108_ _05143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15005_ _02044_ clknet_leaf_375_clk_i memory\[3\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12217_ _06146_ _06422_ _06287_ _06423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_122_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07226__I1 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13197_ _06831_ _02586_ _02588_ _02590_ _02591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_23_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10230__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12148_ _06272_ _06350_ _06352_ _06354_ _06355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06985__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13555__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_10_Right_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12079_ _05686_ _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_159_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_139_Right_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_17_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12435__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15769_ _00728_ clknet_leaf_146_clk_i memory\[62\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_63_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12286__I1 net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08310_ _03948_ _01388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11803__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08384__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09290_ _04214_ memory\[32\]\[15\] _04477_ _04483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_43_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08241_ _03787_ memory\[17\]\[17\] _03904_ _03912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_43_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09279__I _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08172_ _03875_ _01323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12202__A4 _06408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07123_ _03280_ _00869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_319_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07054_ _03242_ _00838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08414__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07217__I1 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10154__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07527__I _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09943__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07956_ _03215_ memory\[19\]\[29\] _03733_ _03743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input28_I data_i[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09914__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06907_ _03135_ memory\[14\]\[3\] _03126_ _03136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11493__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07887_ _03706_ _01207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12674__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_106_Right_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_74_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09626_ _04675_ _01977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07262__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09557_ _04638_ _01945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08508_ _04053_ _01481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_65_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09488_ _04591_ memory\[35\]\[8\] _04575_ _04592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_80_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08439_ _03781_ memory\[20\]\[14\] _04012_ _04017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_22_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_68_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_189_4001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_136_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_4012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11450_ _05660_ _05663_ _05665_ _05666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_191_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_738 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10401_ _05102_ _00245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11381_ _03321_ memory\[62\]\[6\] _05616_ _05623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13120_ _02515_ _00753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07638__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10332_ _03211_ _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10460__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_115_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13051_ _02446_ _02447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10263_ _05017_ _00192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07208__I1 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12002_ _06210_ _06211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_163_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_43_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12901__A2 _02269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10194_ _04591_ memory\[45\]\[8\] _04969_ _04978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10999__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13375__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_121_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07373__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13953_ _00992_ clknet_leaf_326_clk_i memory\[49\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12904_ _03450_ _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07392__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13884_ _00923_ clknet_leaf_283_clk_i memory\[11\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_119_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15623_ _00582_ clknet_leaf_235_clk_i memory\[58\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12835_ _06484_ _02234_ _02235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_268_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15554_ _00513_ clknet_leaf_320_clk_i memory\[56\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12766_ _02165_ _02166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_431_clk_i clknet_5_1__leaf_clk_i clknet_leaf_431_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14505_ _01544_ clknet_leaf_175_clk_i memory\[23\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_12_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12518__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11717_ _05794_ _05930_ _05931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15485_ _00444_ clknet_leaf_333_clk_i memory\[54\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12697_ _06843_ _06862_ _02081_ _02098_ _02099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_72_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11648_ _05767_ _05855_ _05862_ _05863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_14436_ _01475_ clknet_leaf_377_clk_i memory\[21\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput12 data_i[14] net12 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_0_126_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput23 data_i[24] net23 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput34 data_i[5] net34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_320_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07447__I1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14367_ _01406_ clknet_leaf_365_clk_i memory\[1\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11579_ _05661_ _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12454__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07548__S _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10451__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13318_ _02709_ _02710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_14298_ _01337_ clknet_leaf_2_clk_i memory\[29\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_149_24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12579__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13249_ memory\[62\]\[25\] memory\[63\]\[25\] _02448_ _02642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09763__S _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10203__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07810_ _03200_ memory\[6\]\[24\] _03661_ _03666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08790_ _04209_ _01607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_36_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08379__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09562__I _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07741_ _03629_ _01138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_84_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_84_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07672_ _03197_ memory\[10\]\[23\] _03589_ _03593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_9_Left_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07383__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09411_ _04199_ memory\[34\]\[8\] _04538_ _04547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06886__A2 _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09342_ _04510_ _01858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_847 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13081__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09003__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09273_ _04197_ memory\[32\]\[7\] _04466_ _04474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10149__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_62_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08224_ _03770_ memory\[17\]\[9\] _03893_ _03903_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12267__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08155_ _03866_ _01315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07106_ _03271_ _00861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07458__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08086_ _03770_ memory\[15\]\[9\] _03819_ _03829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_101_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_140_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07037_ _03233_ _00830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09673__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_73_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10612__S _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09472__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08988_ _04323_ _01691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07939_ _03734_ _01231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08088__I _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10950_ memory\[55\]\[28\] _03211_ _05385_ _05394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11951__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09609_ _04621_ memory\[36\]\[22\] _04664_ _04667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10881_ _05064_ memory\[54\]\[28\] _05348_ _05357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12620_ _06774_ _06790_ _06805_ _06820_ _06821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__13072__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08816__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07126__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12551_ _06480_ _06752_ _06482_ _06753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__07826__A1 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08874__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_156_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_156_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11502_ _05717_ _05718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_80_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09848__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08752__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15270_ _00229_ clknet_leaf_270_clk_i memory\[47\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12482_ _06639_ _06654_ _06669_ _06684_ _06685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_151_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_117_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14221_ _01260_ clknet_leaf_198_clk_i memory\[12\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11433_ _03373_ memory\[62\]\[31\] _05615_ _05650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_117_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_46_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14152_ _01191_ clknet_leaf_221_clk_i memory\[7\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_134_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11364_ _05613_ _00697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13103_ memory\[30\]\[22\] memory\[31\]\[22\] _02084_ _02499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10315_ _05052_ memory\[46\]\[22\] _05048_ _05053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14083_ _01122_ clknet_leaf_304_clk_i memory\[63\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11295_ _05576_ _00665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07167__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13034_ memory\[30\]\[21\] memory\[31\]\[21\] _02084_ _02431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10246_ _05005_ _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_119_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09051__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10177_ _04968_ _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_156_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14985_ _02024_ clknet_leaf_40_clk_i memory\[38\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_92_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13936_ _00975_ clknet_leaf_124_clk_i memory\[8\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07365__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08927__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13867_ _00906_ clknet_leaf_258_clk_i memory\[39\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11353__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_370_clk_i clknet_5_12__leaf_clk_i clknet_leaf_370_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15606_ _00565_ clknet_leaf_159_clk_i memory\[57\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12818_ memory\[40\]\[18\] memory\[41\]\[18\] memory\[42\]\[18\] memory\[43\]\[18\]
+ _06875_ _02217_ _02218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__13063__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07117__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13798_ _00837_ clknet_leaf_204_clk_i memory\[16\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15537_ _00496_ clknet_leaf_154_clk_i memory\[55\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12248__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12749_ memory\[24\]\[17\] memory\[25\]\[17\] memory\[26\]\[17\] memory\[27\]\[17\]
+ _06472_ _06611_ _02150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08865__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15468_ _00427_ clknet_leaf_275_clk_i memory\[53\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12249__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12692__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_385_clk_i clknet_5_7__leaf_clk_i clknet_leaf_385_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14419_ _01458_ clknet_leaf_99_clk_i memory\[20\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15399_ _00358_ clknet_leaf_293_clk_i memory\[51\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_4_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10424__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07278__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09290__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13118__A2 _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_38_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09960_ _04629_ memory\[41\]\[26\] _04847_ _04854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12912__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08911_ _04243_ memory\[26\]\[29\] _04272_ _04282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_55_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09891_ _04817_ _00020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08842_ _04244_ _01624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10432__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_191_Right_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_323_clk_i clknet_5_10__leaf_clk_i clknet_leaf_323_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12629__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08773_ _04197_ memory\[25\]\[7\] _04183_ _04198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07724_ _03620_ _01130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07356__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07655_ _03172_ memory\[10\]\[15\] _03578_ _03584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11771__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12359__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_338_clk_i clknet_5_9__leaf_clk_i clknet_leaf_338_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11263__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_0_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07586_ _03172_ memory\[0\]\[15\] _03541_ _03547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13054__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09325_ _03305_ net74 _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_138_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_146_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09668__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09256_ _04464_ _01818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08207_ _03894_ _01339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08608__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09187_ _04247_ memory\[30\]\[31\] _04393_ _04428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08138_ _03746_ memory\[29\]\[0\] _03857_ _03858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_151_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_216_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10040__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_75_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08069_ _03820_ _01275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12822__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10100_ _04633_ memory\[43\]\[28\] _04919_ _04928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09033__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11080_ _05058_ memory\[57\]\[25\] _05457_ _05463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12868__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10031_ _04891_ _00086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10342__S _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12332__A3 _06536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output59_I net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14770_ _01809_ clknet_leaf_87_clk_i memory\[31\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11982_ _06191_ _06192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__08747__S _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07651__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13721_ _03340_ memory\[9\]\[15\] _03086_ _03092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10933_ _05362_ _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_158_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_158_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13045__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13652_ _05777_ _03038_ _03039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10864_ _05325_ _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_116_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_17_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12603_ _06318_ _06799_ _06801_ _06803_ _06804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__13140__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08847__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12068__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13583_ _05747_ _02966_ _02968_ _02970_ _02971_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10795_ _05311_ _00430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15322_ _00281_ clknet_leaf_380_clk_i memory\[48\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08482__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12534_ memory\[46\]\[14\] memory\[47\]\[14\] _06596_ _06736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_30_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15253_ _00212_ clknet_leaf_384_clk_i memory\[46\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12465_ _06318_ _06663_ _06665_ _06667_ _06668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10517__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11700__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14204_ _01243_ clknet_leaf_373_clk_i memory\[12\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10406__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11416_ _05641_ _00721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07027__A2 _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12396_ _06325_ _06599_ _06600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15184_ _00143_ clknet_leaf_19_clk_i memory\[44\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14135_ _01174_ clknet_leaf_141_clk_i memory\[6\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11347_ memory\[61\]\[22\] _03193_ _05602_ _05605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09972__A1 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12732__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09024__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14066_ _01105_ clknet_leaf_120_clk_i memory\[10\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12859__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11278_ _03355_ memory\[60\]\[22\] _05565_ _05568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10229_ _04996_ _00179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13017_ memory\[36\]\[21\] memory\[37\]\[21\] _02338_ _02414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07586__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_2_2_0_clk_i clknet_0_clk_i clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_33_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_418_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08657__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14968_ _02007_ clknet_leaf_71_clk_i memory\[37\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07561__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13919_ _00958_ clknet_leaf_309_clk_i memory\[8\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12179__S _06319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14899_ _01938_ clknet_leaf_75_clk_i memory\[35\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07440_ _03468_ _00998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_8_Right_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_165_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07371_ _03166_ memory\[8\]\[13\] _03426_ _03430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08838__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12907__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09110_ _04387_ _01749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09488__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08392__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12890__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09041_ _04237_ memory\[28\]\[26\] _04344_ _04351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09263__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10948__I1 _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13738__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11070__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07736__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09943_ _04612_ memory\[41\]\[18\] _04836_ _04845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_460 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_39_Right_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_262_clk_i clknet_5_24__leaf_clk_i clknet_leaf_262_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10162__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09874_ _04808_ _00012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08825_ _03199_ _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__13473__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13275__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08567__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08756_ _04186_ _01596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input10_I data_i[12] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_277_clk_i clknet_5_13__leaf_clk_i clknet_leaf_277_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07707_ _03611_ _01122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08687_ _03756_ memory\[24\]\[2\] _04146_ _04149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12873__I1 memory\[39\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07638_ _03147_ memory\[10\]\[7\] _03567_ _03575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_48_Right_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_4074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_200_clk_i clknet_5_27__leaf_clk_i clknet_leaf_200_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08829__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07569_ _03147_ memory\[0\]\[7\] _03530_ _03538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11721__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_165_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09308_ _04492_ _01842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10580_ _05197_ _00329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09239_ _04231_ memory\[31\]\[23\] _04452_ _04456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_6_clk_i clknet_5_5__leaf_clk_i clknet_leaf_6_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_181_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11520__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_215_clk_i clknet_5_30__leaf_clk_i clknet_leaf_215_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_185_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12250_ _06453_ _06455_ _06456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_146_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_367_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11201_ _03346_ memory\[5\]\[18\] _05518_ _05527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11061__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12181_ memory\[46\]\[9\] memory\[47\]\[9\] _05907_ _06388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_57_Right_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11132_ _05490_ _00588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__11168__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11063_ _05041_ memory\[57\]\[17\] _05446_ _05454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13502__A2 _02890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11513__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09861__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10014_ _04882_ _00078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14822_ _01861_ clknet_leaf_52_clk_i memory\[33\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07381__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14753_ _01792_ clknet_leaf_412_clk_i memory\[31\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11965_ _06174_ _06175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_157_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_66_Right_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_13704_ _03323_ memory\[9\]\[7\] _03075_ _03083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10875__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_15_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10916_ _05376_ _00486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14684_ _01723_ clknet_leaf_377_clk_i memory\[2\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07740__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11896_ _05741_ _06106_ _06107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13635_ _05719_ _03021_ _05739_ _03022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10847_ _05339_ _00454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13566_ memory\[56\]\[30\] memory\[57\]\[30\] memory\[58\]\[30\] memory\[59\]\[30\]
+ _05711_ _03748_ _02954_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10778_ _05029_ memory\[53\]\[11\] _05301_ _05303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09101__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_915 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15305_ _00264_ clknet_leaf_295_clk_i memory\[48\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12517_ _06717_ _06718_ _06304_ _06719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12526__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13131__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10247__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13497_ _02886_ net60 _02382_ _02887_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15236_ _00195_ clknet_leaf_405_clk_i memory\[46\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08940__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12448_ memory\[8\]\[13\] memory\[9\]\[13\] memory\[10\]\[13\] memory\[11\]\[13\]
+ _06582_ _06032_ _06651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__09245__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_1__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_75_Right_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15167_ _00126_ clknet_leaf_423_clk_i memory\[44\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12379_ memory\[8\]\[12\] memory\[9\]\[12\] memory\[10\]\[12\] memory\[11\]\[12\]
+ _06582_ _06032_ _06583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_188_3987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11752__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14118_ _01157_ clknet_leaf_222_clk_i memory\[6\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15098_ _00057_ clknet_leaf_441_clk_i memory\[41\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11078__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12261__I _03224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06940_ _03160_ memory\[14\]\[11\] _03157_ _03161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_91_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12927__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14049_ _01088_ clknet_leaf_301_clk_i memory\[10\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07559__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I address_i[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11355__I1 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08610_ _03816_ memory\[22\]\[31\] _04072_ _04107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10710__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09590_ _04602_ memory\[36\]\[13\] _04653_ _04657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13257__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_84_Right_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08541_ _04070_ _01497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_385 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08472_ _03814_ memory\[20\]\[30\] _04000_ _04034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07731__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07423_ _03459_ _00990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07354_ _03141_ memory\[8\]\[5\] _03415_ _03421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07285_ _03384_ _00927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09024_ _04220_ memory\[28\]\[18\] _04333_ _04342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_93_Right_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_143_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13468__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11743__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07466__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07411__A2 _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09926_ _04824_ _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_0_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13496__A1 _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07265__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09681__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12838__A4 _02237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09857_ _04799_ _00004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_146_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08808_ _04221_ _01613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08297__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09788_ _04750_ _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_0_Left_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_77_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_107_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08739_ _03808_ memory\[24\]\[27\] _04168_ _04176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11515__I _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11750_ _05724_ _05962_ _05963_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_139_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10701_ _05020_ memory\[52\]\[7\] _05254_ _05262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12547__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11681_ _05724_ _05894_ _05895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_83_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13420_ memory\[30\]\[27\] memory\[31\]\[27\] _05737_ _02811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10632_ _05225_ _00353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11657__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11282__I0 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_154_clk_i clknet_5_18__leaf_clk_i clknet_leaf_154_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10563_ _05188_ _00321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10067__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13351_ memory\[40\]\[26\] memory\[41\]\[26\] memory\[42\]\[26\] memory\[43\]\[26\]
+ _05692_ _02217_ _02743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_36_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09856__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12302_ _06411_ _06499_ _06506_ _06507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_10494_ _05018_ memory\[4\]\[6\] _05145_ _05152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13282_ _02344_ _02674_ _02675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_20_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15021_ _02060_ clknet_leaf_171_clk_i memory\[3\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11034__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12233_ memory\[14\]\[10\] memory\[15\]\[10\] _06302_ _06439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09778__I1 _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_169_clk_i clknet_5_28__leaf_clk_i clknet_leaf_169_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07789__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_113_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12164_ memory\[12\]\[9\] memory\[13\]\[9\] _06025_ _06371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11115_ _05481_ _00580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12909__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12095_ memory\[14\]\[8\] memory\[15\]\[8\] _06302_ _06303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13487__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11046_ _05024_ memory\[57\]\[9\] _05435_ _05445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_183_3895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11593__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11626__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13239__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10530__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14805_ _01844_ clknet_leaf_74_clk_i memory\[32\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08000__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15785_ _00744_ clknet_leaf_260_clk_i net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XFILLER_0_98_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12997_ _06835_ _02393_ _02178_ _02394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_107_clk_i clknet_5_23__leaf_clk_i clknet_leaf_107_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10848__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14736_ _01775_ clknet_leaf_90_clk_i memory\[30\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_8_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08935__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11948_ _06157_ _06158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07713__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12462__A2 _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14667_ _01706_ clknet_leaf_185_clk_i memory\[28\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11879_ _03116_ _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_131_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_38_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11361__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13618_ memory\[16\]\[30\] memory\[17\]\[30\] memory\[18\]\[30\] memory\[19\]\[30\]
+ _05761_ _05762_ _03006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_7_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14598_ _01637_ clknet_leaf_179_clk_i memory\[26\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12845__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13549_ _02501_ _02937_ _02938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_82_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07070_ _03250_ _00846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_41_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09218__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15219_ _00178_ clknet_leaf_14_clk_i memory\[45\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10705__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12073__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07286__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_4__f_clk_i clknet_2_0_0_clk_i clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_10_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13478__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07972_ _03754_ memory\[12\]\[1\] _03752_ _03755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11328__I1 _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09711_ _04587_ memory\[38\]\[6\] _04714_ _04721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06923_ _03147_ memory\[14\]\[7\] _03126_ _03148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13573__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09642_ _04684_ _01984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07952__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_315_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09573_ _04585_ memory\[36\]\[5\] _04642_ _04648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08524_ _03798_ memory\[21\]\[22\] _04059_ _04062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10839__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13650__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07704__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11887__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08455_ _04025_ _01456_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12367__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_102_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07180__I1 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_71_clk_i clknet_5_16__leaf_clk_i clknet_leaf_71_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11271__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07406_ _03218_ memory\[8\]\[30\] _03414_ _03448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_82_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_110_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08386_ _03796_ memory\[1\]\[21\] _03987_ _03989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09457__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13402__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_46_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07337_ _03411_ _00952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09209__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07268_ _03220_ _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_86_clk_i clknet_5_17__leaf_clk_i clknet_leaf_86_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_115_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09007_ _04321_ _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11016__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07199_ _03326_ _00899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_83_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09475__I _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_148_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13181__A3 _02560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13013__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11319__I1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09909_ _04827_ _00028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08196__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_45_Left_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12920_ _02302_ _02309_ _02317_ _02318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10350__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output41_I net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08819__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_24_clk_i clknet_5_4__leaf_clk_i clknet_leaf_24_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12851_ _06835_ _02249_ _02178_ _02250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_122_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_122_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11802_ _05651_ _06005_ _06013_ _06014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_16_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15570_ _00529_ clknet_leaf_164_clk_i memory\[56\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08755__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12782_ _06831_ _02176_ _02179_ _02181_ _02182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_84_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14521_ _01560_ clknet_leaf_106_clk_i memory\[23\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11733_ _05682_ _05945_ _05687_ _05946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_138_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39_clk_i clknet_5_7__leaf_clk_i clknet_leaf_39_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_154_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14452_ _01491_ clknet_leaf_92_clk_i memory\[21\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_25_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11664_ memory\[48\]\[2\] memory\[49\]\[2\] memory\[50\]\[2\] memory\[51\]\[2\] _05692_
+ _05694_ _05878_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_3_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_3_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_54_Left_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13403_ memory\[36\]\[27\] memory\[37\]\[27\] _02338_ _02794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11255__I0 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10615_ _05215_ _00346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14383_ _01422_ clknet_leaf_168_clk_i memory\[1\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08120__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11595_ _05654_ _05805_ _05807_ _05809_ _05810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_107_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11955__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09586__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13334_ memory\[14\]\[26\] memory\[15\]\[26\] _02193_ _02726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08490__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10546_ _05070_ memory\[4\]\[31\] _05144_ _05179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08671__I1 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13265_ _06848_ _02657_ _05791_ _02658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10477_ _05142_ _00281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_185_3924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15004_ _02043_ clknet_leaf_374_clk_i memory\[3\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_264_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12216_ memory\[54\]\[10\] memory\[55\]\[10\] _06421_ _06422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13196_ _06838_ _02589_ _02590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12380__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12147_ _06279_ _06353_ _06354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_63_Left_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07834__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13555__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12078_ memory\[54\]\[8\] memory\[55\]\[8\] _05684_ _06286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_600 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11029_ _05436_ _00539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_86_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13571__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08665__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15768_ _00727_ clknet_leaf_146_clk_i memory\[62\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09687__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_129_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14719_ _01758_ clknet_leaf_412_clk_i memory\[30\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12187__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15699_ _00658_ clknet_leaf_148_clk_i memory\[60\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08240_ _03911_ _01355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_43_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_72_Left_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_129_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09439__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12818__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12199__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08171_ _03785_ memory\[29\]\[16\] _03868_ _03875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11246__I0 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_60_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12915__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07122_ _03156_ memory\[13\]\[10\] _03279_ _03280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07053_ _03160_ memory\[16\]\[11\] _03240_ _03242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10435__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_363 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09611__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13746__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_81_Left_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07744__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07955_ _03742_ _01239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_143_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06906_ _03134_ _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10170__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07886_ _03212_ memory\[7\]\[28\] _03697_ _03706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12674__A2 _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07925__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09625_ _04637_ memory\[36\]\[30\] _04641_ _04675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10685__A1 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13481__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09556_ _04637_ memory\[35\]\[30\] _04574_ _04638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08575__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_90_Left_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08507_ _03781_ memory\[21\]\[14\] _04048_ _04053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09487_ _03149_ _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__08350__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08438_ _04016_ _01448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_22_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12729__A3 _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08369_ _03779_ memory\[1\]\[13\] _03976_ _03980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07919__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10400_ _05060_ memory\[47\]\[26\] _05095_ _05102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11380_ _05622_ _00704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09850__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10331_ _05063_ _00214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13050_ memory\[60\]\[22\] memory\[61\]\[22\] _02164_ _02446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10262_ _05016_ memory\[46\]\[5\] _05006_ _05017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_115_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09602__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12362__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12001_ memory\[60\]\[7\] memory\[61\]\[7\] _05656_ _06210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10193_ _04977_ _00162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_44_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12901__A3 _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_100_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08169__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11176__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13952_ _00991_ clknet_leaf_327_clk_i memory\[49\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_89_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12903_ _02301_ _00750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13883_ _00922_ clknet_leaf_399_clk_i memory\[39\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15622_ _00581_ clknet_leaf_236_clk_i memory\[58\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12834_ memory\[16\]\[18\] memory\[17\]\[18\] memory\[18\]\[18\] memory\[19\]\[18\]
+ _02233_ _06485_ _02234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_115_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15553_ _00512_ clknet_leaf_324_clk_i memory\[56\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12765_ memory\[60\]\[18\] memory\[61\]\[18\] _02164_ _02165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14504_ _01543_ clknet_leaf_175_clk_i memory\[23\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11716_ memory\[16\]\[2\] memory\[17\]\[2\] memory\[18\]\[2\] memory\[19\]\[2\] _05795_
+ _05796_ _05930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_12_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15484_ _00443_ clknet_leaf_332_clk_i memory\[54\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12696_ _06467_ _02090_ _02097_ _02098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_71_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11228__I0 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14435_ _01474_ clknet_leaf_355_clk_i memory\[21\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11647_ _05783_ _05857_ _05859_ _05861_ _05862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_181_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput13 data_i[15] net13 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_142_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput24 data_i[25] net24 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_24_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput35 data_i[6] net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14366_ _01405_ clknet_leaf_364_clk_i memory\[1\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08644__I1 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11578_ _05759_ _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_24_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13317_ memory\[52\]\[26\] memory\[53\]\[26\] _05716_ _02709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10529_ _05170_ _00305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_40_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_172_Right_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14297_ _01336_ clknet_leaf_77_clk_i memory\[29\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13225__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_22__f_clk_i clknet_2_2_0_clk_i clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13248_ _02640_ _02641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_58_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__I0 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13179_ _02367_ _02569_ _02571_ _02573_ _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_20_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07080__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12105__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11086__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07740_ _03197_ memory\[63\]\[23\] _03625_ _03629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_84_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_74_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_84_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07671_ _03592_ _01105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09410_ _04546_ _01890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11814__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13605__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09341_ _04197_ memory\[33\]\[7\] _04502_ _04510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08332__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09272_ _04473_ _01825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08223_ _03902_ _01347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12267__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11919__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_43_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_499 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08154_ _03768_ memory\[29\]\[8\] _03857_ _03866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07105_ _03132_ memory\[13\]\[2\] _03268_ _03271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08085_ _03828_ _01283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07036_ _03135_ memory\[16\]\[3\] _03229_ _03233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09954__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_7_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_179_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07474__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08987_ _04181_ memory\[28\]\[0\] _04322_ _04323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07938_ _03187_ memory\[19\]\[20\] _03733_ _03734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07869_ _03674_ _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_39_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_119_Left_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08571__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_212_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_27_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09608_ _04666_ _01968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10880_ _05356_ _00470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13224__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09539_ _04626_ _01939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11523__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_65_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12550_ memory\[22\]\[14\] memory\[23\]\[14\] _06751_ _06752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_156_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11501_ memory\[12\]\[0\] memory\[13\]\[0\] _05716_ _05717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_156_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12481_ _06467_ _06676_ _06683_ _06684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_149_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10681__I1 _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13455__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14220_ _01259_ clknet_leaf_198_clk_i memory\[12\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07649__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_117_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11432_ _05649_ _00729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_117_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_80_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_128_Left_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_149_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14151_ _01190_ clknet_leaf_245_clk_i memory\[7\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11363_ memory\[61\]\[30\] _03217_ _05579_ _05613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13102_ _05659_ _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_10314_ _03193_ _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14082_ _01121_ clknet_leaf_304_clk_i memory\[63\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11294_ _03371_ memory\[60\]\[30\] _05542_ _05576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13033_ _02429_ _02430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12290__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10245_ _03124_ _04787_ _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__10803__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10176_ net76 _04787_ _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_14984_ _02023_ clknet_leaf_37_clk_i memory\[38\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_137_Left_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13686__I1 net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13935_ _00974_ clknet_leaf_203_clk_i memory\[8\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11634__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11941__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13866_ _00905_ clknet_leaf_258_clk_i memory\[39\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1062 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15605_ _00564_ clknet_leaf_160_clk_i memory\[57\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12817_ _05693_ _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_13797_ _00836_ clknet_leaf_338_clk_i memory\[16\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15536_ _00495_ clknet_leaf_153_clk_i memory\[55\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12748_ _06607_ _02148_ _02086_ _02149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_29_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_691 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10821__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15467_ _00426_ clknet_leaf_296_clk_i memory\[53\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12679_ _06445_ _06870_ _02080_ _02081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XPHY_EDGE_ROW_146_Left_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_25_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12249__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_897 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_414_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07559__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14418_ _01457_ clknet_leaf_99_clk_i memory\[20\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_154_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_128_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__I1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15398_ _00357_ clknet_leaf_293_clk_i memory\[51\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_163_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14349_ _01388_ clknet_leaf_194_clk_i memory\[18\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_40_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_761 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_13_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09774__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13118__A3 _02493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_38_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08910_ _04281_ _01655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_161_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10188__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09890_ _04627_ memory\[40\]\[25\] _04811_ _04817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07294__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07053__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08841_ _04243_ memory\[25\]\[29\] _04225_ _04244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08772_ _03146_ _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_58_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07723_ _03172_ memory\[63\]\[15\] _03614_ _03620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07654_ _03583_ _01097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10360__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09014__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07585_ _03546_ _01065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08305__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09324_ _04500_ _01850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_138_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10112__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08853__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_86_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09255_ _04247_ memory\[31\]\[31\] _04429_ _04464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10663__I1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_106_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08206_ _03746_ memory\[17\]\[0\] _03893_ _03894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09186_ _04427_ _01785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12565__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08137_ _03856_ _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_151_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_151_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07268__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10040__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08068_ _03746_ memory\[15\]\[0\] _03819_ _03820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_101_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_112_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12317__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07019_ net31 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10623__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12868__A2 _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07044__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10030_ _04631_ memory\[42\]\[27\] _04883_ _04891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_430_clk_i clknet_5_1__leaf_clk_i clknet_leaf_430_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08792__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12176__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11981_ memory\[28\]\[6\] memory\[29\]\[6\] _05915_ _06191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13720_ _03091_ _00777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_363_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_445_clk_i clknet_5_1__leaf_clk_i clknet_leaf_445_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10932_ _05384_ _00494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_158_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_158_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13651_ memory\[8\]\[31\] memory\[9\]\[31\] memory\[10\]\[31\] memory\[11\]\[31\]
+ _02473_ _05779_ _03038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10863_ _05347_ _00462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09859__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12602_ _06325_ _06802_ _06803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_155_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13582_ _05759_ _02969_ _02970_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_94_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10794_ _05045_ memory\[53\]\[19\] _05301_ _05311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15321_ _00280_ clknet_leaf_380_clk_i memory\[48\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_109_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12533_ _06734_ _06735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_38_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10654__I1 _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_164_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07379__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15252_ _00211_ clknet_leaf_39_clk_i memory\[46\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12464_ _06325_ _06666_ _06667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_87_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14203_ _01242_ clknet_leaf_398_clk_i memory\[19\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12556__A1 _06703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11415_ _03355_ memory\[62\]\[22\] _05638_ _05641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15183_ _00142_ clknet_leaf_36_clk_i memory\[44\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12395_ memory\[40\]\[12\] memory\[41\]\[12\] memory\[42\]\[12\] memory\[43\]\[12\]
+ _06186_ _06326_ _06599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07027__A3 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09594__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14134_ _01173_ clknet_leaf_141_clk_i memory\[6\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11346_ _05604_ _00688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_1_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09972__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12308__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14065_ _01104_ clknet_leaf_122_clk_i memory\[10\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11277_ _05567_ _00656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13016_ _02319_ _02405_ _02412_ _02413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_10228_ _04625_ memory\[45\]\[24\] _04991_ _04996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08003__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08783__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_33_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_33_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10332__I _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10159_ _04959_ _00146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_50_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14967_ _02006_ clknet_leaf_12_clk_i memory\[37\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07338__I1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13918_ _00957_ clknet_leaf_308_clk_i memory\[8\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10342__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14898_ _01937_ clknet_leaf_76_clk_i memory\[35\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13849_ _00888_ clknet_leaf_109_clk_i memory\[13\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_108_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11163__I _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_18_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07370_ _03429_ _00967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08673__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15519_ _00478_ clknet_leaf_331_clk_i memory\[55\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10708__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12890__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09040_ _04350_ _01716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13339__A3 _02730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_167_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11539__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09942_ _04844_ _00044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10443__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09873_ _04610_ memory\[40\]\[17\] _04800_ _04808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_70_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13754__S _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08824_ _04232_ _01618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10581__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07752__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08755_ _04185_ memory\[25\]\[1\] _04183_ _04186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08526__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11274__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07706_ _03147_ memory\[63\]\[7\] _03603_ _03611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08686_ _04148_ _01564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10333__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07637_ _03574_ _01089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09679__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_192_4064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08583__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07568_ _03537_ _01057_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09307_ _04231_ memory\[32\]\[23\] _04488_ _04492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13502__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_153_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07499_ _03500_ _01025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09478__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09238_ _04455_ _01809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12538__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09169_ _04229_ memory\[30\]\[22\] _04416_ _04419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_131_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_5_31__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07927__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11200_ _05526_ _00620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12180_ _06386_ _06387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_114_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07965__A1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11131_ _03344_ memory\[58\]\[17\] _05482_ _05490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12632__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output71_I net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11062_ _05453_ _00555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13664__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12710__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10013_ _04614_ memory\[42\]\[19\] _04872_ _04882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_129_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08758__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14821_ _01860_ clknet_leaf_402_clk_i memory\[33\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_384_clk_i clknet_5_7__leaf_clk_i clknet_leaf_384_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08517__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14752_ _01791_ clknet_leaf_412_clk_i memory\[31\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11964_ memory\[36\]\[6\] memory\[37\]\[6\] _05733_ _06174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10324__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_1245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13703_ _03082_ _00769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_169_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10915_ memory\[55\]\[11\] _03159_ _05374_ _05376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12079__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14683_ _01722_ clknet_leaf_1_clk_i memory\[28\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11895_ memory\[32\]\[5\] memory\[33\]\[5\] memory\[34\]\[5\] memory\[35\]\[5\] _05742_
+ _05743_ _06106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_15_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_399_clk_i clknet_5_1__leaf_clk_i clknet_leaf_399_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13634_ memory\[54\]\[31\] memory\[55\]\[31\] _05720_ _03021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10846_ _05029_ memory\[54\]\[11\] _05337_ _05339_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10627__I1 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13565_ _05705_ _02952_ _05756_ _02953_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10528__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10777_ _05302_ _00421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15304_ _00263_ clknet_leaf_295_clk_i memory\[48\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12516_ memory\[14\]\[14\] memory\[15\]\[14\] _06302_ _06718_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_322_clk_i clknet_5_10__leaf_clk_i clknet_leaf_322_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13496_ _02840_ _02855_ _02870_ _02885_ _02886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_23_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_670 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15235_ _00194_ clknet_leaf_411_clk_i memory\[46\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12447_ _06028_ _06649_ _06304_ _06650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_2_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_65_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_112_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15166_ _00125_ clknet_leaf_423_clk_i memory\[44\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12378_ _05669_ _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_91_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11359__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_188_3988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14117_ _01156_ clknet_leaf_294_clk_i memory\[6\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_188_3999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_337_clk_i clknet_5_11__leaf_clk_i clknet_leaf_337_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11329_ _05595_ _00680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15097_ _00056_ clknet_leaf_3_clk_i memory\[41\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14048_ _01087_ clknet_leaf_307_clk_i memory\[10\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_34_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10062__I _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_98_1194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08540_ _03814_ memory\[21\]\[30\] _04036_ _04070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10315__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09181__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08471_ _04033_ _01464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_259_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_77_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07422_ memory\[49\]\[3\] _03315_ _03455_ _03459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07353_ _03420_ _00959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07284_ memory\[11\]\[4\] _03317_ _03379_ _03384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_94 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09023_ _04341_ _01708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_311_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08995__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11269__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12379__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09962__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09925_ _04835_ _00036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08747__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13740__I0 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09856_ _04593_ memory\[40\]\[9\] _04789_ _04799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10554__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08807_ _04220_ memory\[25\]\[18\] _04204_ _04221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09787_ _04761_ _02052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06999_ net25 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_107_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08738_ _04175_ _01589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_124_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08669_ memory\[23\]\[26\] _03363_ _04132_ _04139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11732__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10700_ _05261_ _00385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11680_ memory\[8\]\[2\] memory\[9\]\[2\] memory\[10\]\[2\] memory\[11\]\[2\] _05893_
+ _05726_ _05894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_48_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_120_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12759__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13232__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10631_ memory\[51\]\[6\] _03143_ _05218_ _05225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12627__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10348__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_113_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13350_ _02213_ _02741_ _02352_ _02742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_106_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_631 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10562_ _05018_ memory\[50\]\[6\] _05181_ _05188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_573 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_45_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12301_ _06142_ _06501_ _06503_ _06505_ _06506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_17_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13281_ memory\[32\]\[25\] memory\[33\]\[25\] memory\[34\]\[25\] memory\[35\]\[25\]
+ _02205_ _02345_ _02674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_10493_ _05151_ _00288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_101_Left_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07657__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15020_ _02059_ clknet_leaf_169_clk_i memory\[3\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12232_ _06437_ _06438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_20_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11687__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08840__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12163_ _06155_ _06365_ _06367_ _06369_ _06370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_11114_ _03327_ memory\[58\]\[9\] _05471_ _05481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_9_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12094_ _05683_ _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_9_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11045_ _05444_ _00547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11498__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08488__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10811__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07392__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11593__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_99_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14804_ _01843_ clknet_leaf_76_clk_i memory\[32\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07191__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12996_ memory\[54\]\[21\] memory\[55\]\[21\] _02312_ _02393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15784_ _00743_ clknet_leaf_260_clk_i net43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_86_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14735_ _01774_ clknet_leaf_127_clk_i memory\[30\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11947_ memory\[4\]\[6\] memory\[5\]\[6\] _06156_ _06157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_260_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14666_ _01705_ clknet_leaf_183_clk_i memory\[28\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11878_ _05705_ _06088_ _06018_ _06089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_86_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13617_ _05753_ _03004_ _05687_ _03005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_157_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10829_ _05012_ memory\[54\]\[3\] _05326_ _05330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14597_ _01636_ clknet_leaf_408_clk_i memory\[26\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_261_clk_i clknet_5_24__leaf_clk_i clknet_leaf_261_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_6_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12845__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13548_ memory\[24\]\[29\] memory\[25\]\[29\] memory\[26\]\[29\] memory\[27\]\[29\]
+ _02363_ _02502_ _02937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_55_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13569__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13479_ _05676_ _02864_ _02866_ _02868_ _02869_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_129_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07567__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15218_ _00177_ clknet_leaf_14_clk_i memory\[45\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07229__I0 memory\[39\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_276_clk_i clknet_5_12__leaf_clk_i clknet_leaf_276_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_140_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08977__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15149_ _00108_ clknet_leaf_24_clk_i memory\[43\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10784__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09782__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07971_ _03128_ _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08729__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13478__A2 _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09710_ _04720_ _02016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11817__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06922_ _03146_ _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08398__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10536__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09641_ _04585_ memory\[37\]\[5\] _04678_ _04684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_5_clk_i clknet_5_4__leaf_clk_i clknet_leaf_5_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_136_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_214_clk_i clknet_5_30__leaf_clk_i clknet_leaf_214_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09572_ _04647_ _01951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09154__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08523_ _04061_ _01488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_141_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08901__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08454_ _03796_ memory\[20\]\[21\] _04023_ _04025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_65_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09022__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07405_ _03447_ _00984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_186_Right_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_148_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_229_clk_i clknet_5_26__leaf_clk_i clknet_leaf_229_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08385_ _03988_ _01423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10168__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_82_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07336_ memory\[11\]\[29\] _03369_ _03401_ _03411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08861__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07267_ _03372_ _00921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12383__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09006_ _04332_ _01700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07198_ memory\[39\]\[8\] _03325_ _03309_ _03326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07640__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13013__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_6_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13713__I0 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09908_ _04577_ memory\[41\]\[1\] _04825_ _04827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10631__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09839_ _04790_ _02075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13227__B _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12772__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08101__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_161_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_161_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11526__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12850_ memory\[54\]\[19\] memory\[55\]\[19\] _06421_ _02249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07940__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_122_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11801_ _05676_ _06007_ _06009_ _06012_ _06013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_90_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12781_ _06838_ _02180_ _02181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_96_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14520_ _01559_ clknet_leaf_108_clk_i memory\[23\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_95_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11732_ memory\[54\]\[3\] memory\[55\]\[3\] _05684_ _05945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_90_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_138_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14451_ _01490_ clknet_leaf_99_clk_i memory\[21\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11663_ _05682_ _05876_ _05687_ _05877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_166_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_153_Right_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_25_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_25_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13402_ _02319_ _02785_ _02792_ _02793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_10614_ _05070_ memory\[50\]\[31\] _05180_ _05215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09867__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14382_ _01421_ clknet_leaf_169_clk_i memory\[1\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11594_ _05668_ _05808_ _05809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_49_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13333_ _02724_ _02725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_107_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10545_ _05178_ _00313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_107_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13264_ memory\[6\]\[25\] memory\[7\]\[25\] _02322_ _02657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10476_ _05068_ memory\[48\]\[30\] _05108_ _05142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_207_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12306__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15003_ _02042_ clknet_leaf_399_clk_i memory\[38\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_62_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12215_ _05683_ _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_185_3925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13195_ memory\[48\]\[24\] memory\[49\]\[24\] memory\[50\]\[24\] memory\[51\]\[24\]
+ _05725_ _06839_ _02589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_138_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12146_ memory\[56\]\[9\] memory\[57\]\[9\] memory\[58\]\[9\] memory\[59\]\[9\] _06138_
+ _06280_ _06353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_124_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13704__I0 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12077_ _06284_ _06285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_159_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09107__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11028_ _05004_ memory\[57\]\[0\] _05435_ _05436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11191__I0 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12041__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_86_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08946__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12976__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12979_ memory\[16\]\[20\] memory\[17\]\[20\] memory\[18\]\[20\] memory\[19\]\[20\]
+ _02233_ _02376_ _02377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15767_ _00726_ clknet_leaf_150_clk_i memory\[62\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09836__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14718_ _01757_ clknet_leaf_414_clk_i memory\[30\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07698__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15698_ _00657_ clknet_leaf_147_clk_i memory\[60\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_129_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14649_ _01688_ clknet_leaf_79_clk_i memory\[27\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_120_Right_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12818__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08170_ _03874_ _01322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13299__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07121_ _03267_ _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_27_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10716__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13148__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07297__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07052_ _03241_ _00837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_43 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07870__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13098__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07096__I _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07954_ _03212_ memory\[19\]\[28\] _03733_ _03742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10451__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10509__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09375__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13320__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06905_ net32 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_143_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07885_ _03705_ _01206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_153_clk_i clknet_5_18__leaf_clk_i clknet_leaf_153_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_409_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11182__I0 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09624_ _04674_ _01976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11882__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10685__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09127__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07760__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11790__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09555_ _03217_ _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_167_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11282__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08506_ _04052_ _01480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_77_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_168_clk_i clknet_5_25__leaf_clk_i clknet_leaf_168_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09486_ _04590_ _01922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_3_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_862 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_849 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_156_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08437_ _03779_ memory\[20\]\[13\] _04012_ _04016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_22_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09687__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13387__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08368_ _03979_ _01415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_34_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_4014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07319_ _03402_ _00943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12985__I1 net52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08299_ _03777_ memory\[18\]\[12\] _03940_ _03943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13002__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13139__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10330_ _05062_ memory\[46\]\[27\] _05048_ _05063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07861__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12126__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_167_3600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10261_ _03140_ _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_115_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12841__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_106_clk_i clknet_5_21__leaf_clk_i clknet_leaf_106_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12000_ _06209_ _00737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07935__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07613__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10192_ _04589_ memory\[45\]\[7\] _04969_ _04977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12901__A4 _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_163_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_895 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_180_3833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09366__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13951_ _00990_ clknet_leaf_347_clk_i memory\[49\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13672__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12902_ _02300_ net50 _06491_ _02301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11873__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13882_ _00921_ clknet_leaf_27_clk_i memory\[39\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07670__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12796__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_159_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12833_ _05691_ _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15621_ _00580_ clknet_leaf_318_clk_i memory\[58\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12288__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13170__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11625__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12764_ _05655_ _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15552_ _00511_ clknet_leaf_324_clk_i memory\[56\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14503_ _01542_ clknet_leaf_172_clk_i memory\[23\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11715_ _05788_ _05928_ _05792_ _05929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_56_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15483_ _00442_ clknet_leaf_374_clk_i memory\[53\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12695_ _06476_ _02092_ _02094_ _02096_ _02097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_51_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13378__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14434_ _01473_ clknet_leaf_358_clk_i memory\[21\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11646_ _05794_ _05860_ _05861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_108_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput14 data_i[16] net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_0_64_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput25 data_i[26] net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14365_ _01404_ clknet_leaf_375_clk_i memory\[1\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10536__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput36 data_i[7] net36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11577_ _05788_ _05790_ _05792_ _05793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10987__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13316_ _02163_ _02703_ _02705_ _02707_ _02708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_161_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10528_ _05052_ memory\[4\]\[22\] _05167_ _05170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08006__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14296_ _01335_ clknet_leaf_85_clk_i memory\[29\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_358_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13225__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13247_ memory\[60\]\[25\] memory\[61\]\[25\] _02164_ _02640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10335__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10459_ _05133_ _00272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10739__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13550__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13178_ _02375_ _02572_ _02573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10271__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12129_ _05914_ _06332_ _06334_ _06336_ _06337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_70_clk_i clknet_5_16__leaf_clk_i clknet_leaf_70_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07644__I _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13302__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_410_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11164__I0 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_84_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07670_ _03194_ memory\[10\]\[22\] _03589_ _03592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09109__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07580__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_85_clk_i clknet_5_17__leaf_clk_i clknet_leaf_85_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15819_ _00778_ clknet_leaf_209_clk_i memory\[9\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09340_ _04509_ _01857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11616__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13081__A3 _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09271_ _04195_ memory\[32\]\[6\] _04466_ _04473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13369__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08222_ _03768_ memory\[17\]\[8\] _03893_ _03902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12041__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08153_ _03865_ _01314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_99_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10978__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09832__I1 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07104_ _03270_ _00860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_23_clk_i clknet_5_5__leaf_clk_i clknet_leaf_23_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_67_1074 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08084_ _03768_ memory\[15\]\[8\] _03819_ _03828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07035_ _03232_ _00829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_77_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09596__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_41_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13541__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_38_clk_i clknet_5_7__leaf_clk_i clknet_leaf_38_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_82_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08986_ _04321_ _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_input33_I data_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09970__S _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07554__I _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09348__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07937_ _03710_ _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11855__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07868_ _03696_ _01198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07490__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09607_ _04619_ memory\[36\]\[21\] _04664_ _04666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07799_ _03184_ memory\[6\]\[19\] _03650_ _03660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11607__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09538_ _04625_ memory\[35\]\[24\] _04617_ _04626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09469_ _03131_ _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_54_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11740__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11500_ _05677_ _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_156_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12480_ _06476_ _06678_ _06680_ _06682_ _06683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_156_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13455__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11431_ _03371_ memory\[62\]\[30\] _05615_ _05649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10356__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12635__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_117_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_565 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14150_ _01189_ clknet_leaf_222_clk_i memory\[7\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_61_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07834__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11362_ _05612_ _00696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_134_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_81_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13101_ _02496_ _02497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_85_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10313_ _05051_ _00208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14081_ _01120_ clknet_leaf_305_clk_i memory\[63\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11293_ _05575_ _00664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_131_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13032_ memory\[28\]\[21\] memory\[29\]\[21\] _06604_ _02429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12966__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11695__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10244_ _03110_ _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11394__I0 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11187__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10175_ _04967_ _00154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09339__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09880__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12099__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11146__I0 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14983_ _02022_ clknet_leaf_40_clk_i memory\[38\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11915__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13934_ _00973_ clknet_leaf_214_clk_i memory\[8\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11846__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08496__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_88_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11941__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13865_ _00904_ clknet_leaf_267_clk_i memory\[39\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15604_ _00563_ clknet_leaf_166_clk_i memory\[57\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12816_ _05689_ _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_13796_ _00835_ clknet_leaf_368_clk_i memory\[16\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_186_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15535_ _00494_ clknet_leaf_241_clk_i memory\[55\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12747_ memory\[30\]\[17\] memory\[31\]\[17\] _02084_ _02148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11650__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10821__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12678_ _06318_ _06872_ _06874_ _06877_ _02080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_15466_ _00425_ clknet_leaf_296_clk_i memory\[53\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_13_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14417_ _01456_ clknet_leaf_100_clk_i memory\[20\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11629_ _05753_ _05843_ _05757_ _05844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08078__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15397_ _00356_ clknet_leaf_313_clk_i memory\[51\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09814__I1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14348_ _01387_ clknet_leaf_193_clk_i memory\[18\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13577__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14279_ _01318_ clknet_leaf_176_clk_i memory\[29\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_104_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11385__I0 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_55_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08840_ _03214_ _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__08250__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08771_ _04196_ _01601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11825__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07722_ _03619_ _01129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_135_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06919__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07653_ _03169_ memory\[10\]\[14\] _03578_ _03583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07584_ _03169_ memory\[0\]\[14\] _03541_ _03546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09323_ _04247_ memory\[32\]\[31\] _04465_ _04500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_138_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_138_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11696__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_29_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09254_ _04463_ _01817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08205_ _03892_ _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12014__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09185_ _04245_ memory\[30\]\[30\] _04393_ _04427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09805__I1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_21__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07816__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08136_ net76 _03855_ _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_43_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_151_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07292__I1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08067_ _03818_ _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_114_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10904__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_112_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09569__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07018_ _03219_ _00825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12948__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08241__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08969_ _04233_ memory\[27\]\[24\] _04308_ _04313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12176__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11980_ _05731_ _06181_ _06189_ _06190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__09741__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09205__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_306_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10931_ memory\[55\]\[19\] _03183_ _05374_ _05384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_158_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13125__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13650_ _05772_ _03036_ _05775_ _03037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10862_ _05045_ memory\[54\]\[19\] _05337_ _05347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_66_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12601_ memory\[40\]\[15\] memory\[41\]\[15\] memory\[42\]\[15\] memory\[43\]\[15\]
+ _06186_ _06326_ _06802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_175_3743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13581_ memory\[0\]\[30\] memory\[1\]\[30\] memory\[2\]\[30\] memory\[3\]\[30\] _05784_
+ _03226_ _02969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_155_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10793_ _05310_ _00429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12566__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12532_ memory\[44\]\[14\] memory\[45\]\[14\] _06319_ _06734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15320_ _00279_ clknet_leaf_380_clk_i memory\[48\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08843__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_109_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_87_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12463_ memory\[40\]\[13\] memory\[41\]\[13\] memory\[42\]\[13\] memory\[43\]\[13\]
+ _06186_ _06326_ _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__10086__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15251_ _00210_ clknet_leaf_40_clk_i memory\[46\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_10_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11414_ _05640_ _00720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14202_ _01241_ clknet_leaf_28_clk_i memory\[19\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09875__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12556__A2 _06725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15182_ _00141_ clknet_leaf_34_clk_i memory\[44\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12394_ _06322_ _06597_ _06461_ _06598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_22_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13397__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14133_ _01172_ clknet_leaf_137_clk_i memory\[6\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11345_ memory\[61\]\[21\] _03190_ _05602_ _05604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08480__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13505__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14064_ _01103_ clknet_leaf_123_clk_i memory\[10\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11276_ _03353_ memory\[60\]\[21\] _05565_ _05567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13015_ _06713_ _02407_ _02409_ _02411_ _02412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10227_ _04995_ _00178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07194__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09980__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_33_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10158_ _04623_ memory\[44\]\[23\] _04955_ _04959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11119__I0 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_50_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_2_3_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10089_ _04922_ _00113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14966_ _02005_ clknet_leaf_13_clk_i memory\[37\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09115__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09732__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13917_ _00956_ clknet_leaf_287_clk_i memory\[8\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12492__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11444__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14897_ _01936_ clknet_leaf_69_clk_i memory\[35\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_18_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08954__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13848_ _00887_ clknet_leaf_138_clk_i memory\[13\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08299__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12476__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13779_ _00818_ clknet_leaf_120_clk_i memory\[14\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_30_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_17_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15518_ _00477_ clknet_leaf_332_clk_i memory\[55\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_31_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_5_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15449_ _00408_ clknet_leaf_269_clk_i memory\[52\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_44_159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_57_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10724__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13100__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_255_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09941_ _04610_ memory\[41\]\[17\] _04836_ _04844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10523__I _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09872_ _04807_ _00011_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_70_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10030__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08823_ _04231_ memory\[25\]\[23\] _04225_ _04232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08754_ _03128_ _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_139_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07705_ _03610_ _01121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08685_ _03754_ memory\[24\]\[1\] _04146_ _04148_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_178_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13107__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07636_ _03144_ memory\[10\]\[6\] _03567_ _03574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_192_4065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07567_ _03144_ memory\[0\]\[6\] _03530_ _03537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11290__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09306_ _04491_ _01841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07498_ memory\[59\]\[6\] _03321_ _03493_ _03500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09237_ _04229_ memory\[31\]\[22\] _04452_ _04455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_146_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_479 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09695__S _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09168_ _04418_ _01776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_131_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_131_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08119_ _03846_ _01299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08462__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09099_ _04227_ memory\[2\]\[21\] _04380_ _04382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_165_Left_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_43_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09494__I _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11130_ _05489_ _00587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07965__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11061_ _05039_ memory\[57\]\[16\] _05446_ _05453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08214__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output64_I net64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10012_ _04881_ _00077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09962__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14820_ _01859_ clknet_leaf_401_clk_i memory\[33\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_4_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14751_ _01790_ clknet_leaf_411_clk_i memory\[31\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11963_ _05699_ _06165_ _06172_ _06173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_98_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_174_Left_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_86_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13702_ _03321_ memory\[9\]\[6\] _03075_ _03082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10914_ _05375_ _00485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11894_ _05736_ _06104_ _05739_ _06105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_58_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14682_ _01721_ clknet_leaf_2_clk_i memory\[28\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13633_ _03019_ _03020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10845_ _05338_ _00453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10809__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10088__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13564_ memory\[62\]\[30\] memory\[63\]\[30\] _02448_ _02952_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10776_ _05026_ memory\[53\]\[10\] _05301_ _05302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15303_ _00262_ clknet_leaf_295_clk_i memory\[48\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12515_ _05681_ _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_136_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13495_ _02358_ _02877_ _02884_ _02885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_48_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_12446_ memory\[14\]\[13\] memory\[15\]\[13\] _06302_ _06649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15234_ _00193_ clknet_leaf_404_clk_i memory\[46\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_23_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_183_Left_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12377_ _06028_ _06580_ _06304_ _06581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15165_ _00124_ clknet_leaf_425_clk_i memory\[44\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10544__S _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_91_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14116_ _01155_ clknet_leaf_294_clk_i memory\[6\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11328_ memory\[61\]\[13\] _03165_ _05591_ _05595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_188_3989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15096_ _00055_ clknet_leaf_7_clk_i memory\[41\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11439__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_52_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14047_ _01086_ clknet_leaf_285_clk_i memory\[10\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11259_ _03336_ memory\[60\]\[13\] _05554_ _05558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07853__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11375__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_192_Left_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_167_Right_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_167_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09705__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14949_ _01988_ clknet_leaf_431_clk_i memory\[37\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12465__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_49_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08470_ _03812_ memory\[20\]\[29\] _04023_ _04033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07421_ _03458_ _00989_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12217__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10079__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07352_ _03138_ memory\[8\]\[4\] _03415_ _03420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07283_ _03383_ _00926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09022_ _04218_ memory\[28\]\[17\] _04333_ _04341_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_14_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_444_clk_i clknet_5_4__leaf_clk_i clknet_leaf_444_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07827__I _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12379__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09924_ _04593_ memory\[41\]\[9\] _04825_ _04835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08859__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12889__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10003__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13496__A3 _02870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11793__B _06002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09855_ _04798_ _00003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_146_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_146_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08806_ _03180_ _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06998_ _03204_ _00820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09786_ memory\[3\]\[9\] _03152_ _04751_ _04761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08737_ _03806_ memory\[24\]\[26\] _04168_ _04175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_134_Right_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_1_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08594__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08668_ _04138_ _01556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07619_ _03221_ memory\[0\]\[31\] _03529_ _03564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08599_ _04101_ _01524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10629__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11812__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10630_ _05224_ _00352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06906__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10561_ _05187_ _00320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07486__I1 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08683__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_392 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12300_ _06149_ _06504_ _06505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07938__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10490__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13280_ _02341_ _02672_ _06866_ _02673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10492_ _05016_ memory\[4\]\[5\] _05145_ _05151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11968__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12231_ memory\[12\]\[10\] memory\[13\]\[10\] _06025_ _06437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08435__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_20_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10364__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10242__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12162_ _06162_ _06368_ _06369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_130_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06997__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11113_ _05480_ _00579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12093_ _06300_ _06301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_TAPCELL_ROW_9_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11044_ _05022_ memory\[57\]\[8\] _05435_ _05444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09935__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_183_3886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_183_3897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11195__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14803_ _01842_ clknet_leaf_79_clk_i memory\[32\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12447__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15783_ _00742_ clknet_leaf_253_clk_i net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XPHY_EDGE_ROW_101_Right_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12995_ _02391_ _02392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_54_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_58_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14734_ _01773_ clknet_leaf_131_clk_i memory\[30\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_203_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11946_ _05701_ _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_169_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14665_ _01704_ clknet_leaf_181_clk_i memory\[28\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11877_ memory\[6\]\[5\] memory\[7\]\[5\] _05706_ _06088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13616_ memory\[22\]\[30\] memory\[23\]\[30\] _05754_ _03004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_16__f_clk_i clknet_2_2_0_clk_i clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10828_ _05329_ _00445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08009__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14596_ _01635_ clknet_leaf_406_clk_i memory\[26\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10338__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12754__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13547_ _02498_ _02935_ _05665_ _02936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10759_ _05010_ memory\[53\]\[2\] _05290_ _05293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_152_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11878__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13478_ _05690_ _02867_ _02868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_15217_ _00176_ clknet_leaf_15_clk_i memory\[45\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10274__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08426__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12429_ memory\[52\]\[13\] memory\[53\]\[13\] _06143_ _06632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07229__I1 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15148_ _00107_ clknet_leaf_24_clk_i memory\[43\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_11_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07970_ _03753_ _01243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08679__S _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15079_ _00038_ clknet_leaf_22_clk_i memory\[41\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06921_ net36 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_93_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09640_ _04683_ _01983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09571_ _04583_ memory\[36\]\[4\] _04642_ _04647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08522_ _03796_ memory\[21\]\[21\] _04059_ _04061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11833__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_95 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_141_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07165__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06927__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09303__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08453_ _04024_ _01455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_65_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_368 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10449__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_102_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07404_ _03215_ memory\[8\]\[29\] _03437_ _03447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_722 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08384_ _03793_ memory\[1\]\[20\] _03987_ _03988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_129_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13402__A3 _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07335_ _03410_ _00951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12610__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07468__I1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_34_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_405_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10472__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07266_ memory\[39\]\[30\] _03371_ _03308_ _03372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_383_clk_i clknet_5_7__leaf_clk_i clknet_leaf_383_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09005_ _04201_ memory\[28\]\[9\] _04322_ _04332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_61_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10184__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07197_ _03149_ _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10224__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_152_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_398_clk_i clknet_5_6__leaf_clk_i clknet_leaf_398_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_6_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09907_ _04826_ _00027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12677__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12772__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09838_ _04573_ memory\[40\]\[0\] _04789_ _04790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_161_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_321_clk_i clknet_5_10__leaf_clk_i clknet_leaf_321_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_38_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12839__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09769_ _04752_ _02043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11800_ _05690_ _06011_ _06012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_69_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12780_ memory\[48\]\[18\] memory\[49\]\[18\] memory\[50\]\[18\] memory\[51\]\[18\]
+ _06699_ _06839_ _02180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_11731_ _05943_ _05944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_90_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12638__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_336_clk_i clknet_5_8__leaf_clk_i clknet_leaf_336_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__06903__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14450_ _01489_ clknet_leaf_98_clk_i memory\[21\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11662_ memory\[54\]\[2\] memory\[55\]\[2\] _05684_ _05876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_25_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_14_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13401_ _05768_ _02787_ _02789_ _02791_ _02792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_107_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_77_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10613_ _05214_ _00345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14381_ _01420_ clknet_leaf_171_clk_i memory\[1\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11593_ memory\[56\]\[1\] memory\[57\]\[1\] memory\[58\]\[1\] memory\[59\]\[1\] _05670_
+ _05671_ _05808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_37_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12574__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07668__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09947__I _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13332_ memory\[12\]\[26\] memory\[13\]\[26\] _05769_ _02724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10544_ _05068_ memory\[4\]\[30\] _05144_ _05178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10094__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13157__A2 _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13263_ _02655_ _02656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10475_ _05141_ _00280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15002_ _02041_ clknet_leaf_430_clk_i memory\[38\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10215__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12214_ _06419_ _06420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_161_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13194_ _06835_ _02587_ _02178_ _02588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_185_3926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12145_ _06276_ _06351_ _06001_ _06352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08499__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09908__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12076_ memory\[52\]\[8\] memory\[53\]\[8\] _06143_ _06284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11027_ _05434_ _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_159_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15835_ _00794_ clknet_leaf_387_clk_i memory\[9\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_354_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15766_ _00725_ clknet_leaf_150_clk_i memory\[62\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07147__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12978_ _05693_ _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_133_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09836__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09123__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14717_ _01756_ clknet_leaf_391_clk_i memory\[30\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08895__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11929_ memory\[56\]\[6\] memory\[57\]\[6\] memory\[58\]\[6\] memory\[59\]\[6\] _06138_
+ _05671_ _06139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15697_ _00656_ clknet_leaf_162_clk_i memory\[60\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_131_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11452__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14648_ _01687_ clknet_leaf_77_clk_i memory\[27\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_429 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_7_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14579_ _01618_ clknet_leaf_95_clk_i memory\[25\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_60_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07578__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_60_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07120_ _03278_ _00868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07051_ _03156_ memory\[16\]\[10\] _03240_ _03241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09793__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11828__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07953_ _03741_ _01238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13328__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08202__S _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06904_ _03133_ _00797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_103_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07884_ _03209_ memory\[7\]\[27\] _03697_ _03705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07386__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09623_ _04635_ memory\[36\]\[29\] _04664_ _04674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09554_ _04636_ _01944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07138__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09033__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08505_ _03779_ memory\[21\]\[13\] _04048_ _04052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08886__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09485_ _04589_ memory\[35\]\[7\] _04575_ _04590_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10693__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09968__S _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08436_ _04015_ _01447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08872__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08367_ _03777_ memory\[1\]\[12\] _03976_ _03979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_68_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_4015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09767__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07318_ memory\[11\]\[20\] _03350_ _03401_ _03402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07488__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10445__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08298_ _03942_ _01382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_119_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13139__A2 _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_132_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07249_ _03360_ _00915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10260_ _05015_ _00191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09063__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__14695__CLK clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11738__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08810__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12921__I _03114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10191_ _04976_ _00161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10642__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_163_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08112__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13698__I0 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11537__I _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_260_clk_i clknet_5_24__leaf_clk_i clknet_leaf_260_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_180_3845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13950_ _00989_ clknet_leaf_347_clk_i memory\[49\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07377__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09007__I _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12901_ _02254_ _02269_ _02284_ _02299_ _02300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_0_92_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13881_ _00920_ clknet_leaf_66_clk_i memory\[39\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_193_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15620_ _00579_ clknet_leaf_318_clk_i memory\[58\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12832_ _06480_ _02231_ _06482_ _02232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08846__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_275_clk_i clknet_5_13__leaf_clk_i clknet_leaf_275_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_139_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15551_ _00510_ clknet_leaf_326_clk_i memory\[56\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_179_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13170__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12763_ _05653_ _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_57_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_178_3796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14502_ _01541_ clknet_leaf_172_clk_i memory\[23\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11714_ memory\[22\]\[2\] memory\[23\]\[2\] _05789_ _05928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15482_ _00441_ clknet_leaf_380_clk_i memory\[53\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12694_ _06484_ _02095_ _02096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_84_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14433_ _01472_ clknet_leaf_353_clk_i memory\[21\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_9 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11645_ memory\[16\]\[1\] memory\[17\]\[1\] memory\[18\]\[1\] memory\[19\]\[1\] _05795_
+ _05796_ _05860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_65_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10817__S _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07398__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput15 data_i[17] net15 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14364_ _01403_ clknet_leaf_374_clk_i memory\[1\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput26 data_i[27] net26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_11576_ _05791_ _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xinput37 data_i[8] net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_0_134_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13315_ _02170_ _02706_ _02707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_24_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10527_ _05169_ _00304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_4_clk_i clknet_5_4__leaf_clk_i clknet_leaf_4_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_150_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14295_ _01334_ clknet_leaf_85_clk_i memory\[29\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07197__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_213_clk_i clknet_5_30__leaf_clk_i clknet_leaf_213_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_122_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13246_ _02639_ _00755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10458_ _05050_ memory\[48\]\[21\] _05131_ _05133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12889__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12433__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08801__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10552__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13177_ memory\[16\]\[23\] memory\[17\]\[23\] memory\[18\]\[23\] memory\[19\]\[23\]
+ _02233_ _02376_ _02572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10389_ _05096_ _00239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12128_ _05921_ _06335_ _06336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_228_clk_i clknet_5_26__leaf_clk_i clknet_leaf_228_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_97_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12059_ _05783_ _06263_ _06265_ _06267_ _06268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07861__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11383__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_31__f_clk_i clknet_2_3_0_clk_i clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15818_ _00777_ clknet_leaf_210_clk_i memory\[9\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12278__I _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15749_ _00708_ clknet_leaf_303_clk_i memory\[62\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11616__A2 _05830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_100_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09270_ _04472_ _01824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_502 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08221_ _03901_ _01346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_23_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_8_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_145_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13103__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08152_ _03766_ memory\[29\]\[7\] _03857_ _03865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_11__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_99_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12227__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07101__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07103_ _03129_ memory\[13\]\[1\] _03268_ _03270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08083_ _03827_ _01282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07034_ _03132_ memory\[16\]\[2\] _03229_ _03232_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09045__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06940__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_796 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_77_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11558__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10462__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_474 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_25_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08985_ _03750_ _03855_ _04321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__10261__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07936_ _03732_ _01230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08867__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input26_I data_i[27] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07867_ _03184_ memory\[7\]\[19\] _03686_ _03696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10902__I1 _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09606_ _04665_ _01967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13057__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07798_ _03659_ _01165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_27_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09537_ _03199_ _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08859__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11607__A2 _05821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12804__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_182_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09468_ _04578_ _01916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08419_ _04006_ _01439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_175_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_156_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10637__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11820__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09399_ _04187_ memory\[34\]\[2\] _04538_ _04541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09497__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10418__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11430_ _05648_ _00728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08107__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06914__I _03140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09284__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11361_ memory\[61\]\[29\] _03214_ _05602_ _05612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_421 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_302_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07946__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13100_ memory\[28\]\[22\] memory\[29\]\[22\] _02495_ _02496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10312_ _05050_ memory\[46\]\[21\] _05048_ _05051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14080_ _01119_ clknet_leaf_306_clk_i memory\[63\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11292_ _03369_ memory\[60\]\[29\] _05565_ _05575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12415__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12651__I _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10243_ _05003_ _00186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13031_ _02336_ _02420_ _02427_ _02428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__12966__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10174_ _04639_ memory\[44\]\[31\] _04932_ _04967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14982_ _02021_ clknet_leaf_40_clk_i memory\[38\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13933_ _00972_ clknet_leaf_209_clk_i memory\[8\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12600__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13864_ _00903_ clknet_leaf_272_clk_i memory\[39\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07770__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15603_ _00562_ clknet_leaf_165_clk_i memory\[57\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12815_ _02213_ _02214_ _06461_ _02215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_186_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13795_ _00834_ clknet_leaf_341_clk_i memory\[16\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_186_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15534_ _00493_ clknet_leaf_257_clk_i memory\[55\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12746_ _02146_ _02147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_57_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09401__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_166_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15465_ _00424_ clknet_leaf_296_clk_i memory\[53\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12677_ _06325_ _06876_ _06877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_5_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14416_ _01455_ clknet_leaf_100_clk_i memory\[20\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_831 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11628_ memory\[46\]\[1\] memory\[47\]\[1\] _05754_ _05843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09275__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15396_ _00355_ clknet_leaf_313_clk_i memory\[51\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_771 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_152_clk_i clknet_5_19__leaf_clk_i clknet_leaf_152_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11082__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14347_ _01386_ clknet_leaf_194_clk_i memory\[18\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11559_ _05664_ _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_123_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11782__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11886__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14278_ _01317_ clknet_leaf_179_clk_i memory\[29\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13229_ memory\[28\]\[24\] memory\[29\]\[24\] _02495_ _02623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_55_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_199_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08770_ _04195_ memory\[25\]\[6\] _04183_ _04196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_72_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_85_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_97_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08687__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07721_ _03169_ memory\[63\]\[14\] _03614_ _03619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_69_Left_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07652_ _03582_ _01096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07583_ _03545_ _01064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_251_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_105_clk_i clknet_5_21__leaf_clk_i clknet_leaf_105_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11841__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09322_ _04499_ _01849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_138_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11696__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09311__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09253_ _04245_ memory\[31\]\[30\] _04429_ _04463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_12_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08204_ _03225_ net75 _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_69_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09184_ _04426_ _01784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13211__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08135_ _03854_ _03855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_78_Left_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_151_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11773__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07766__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09018__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08066_ _03115_ _03306_ _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_102_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07017_ _03218_ memory\[14\]\[30\] _03125_ _03219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_112_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_113_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11288__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10192__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12948__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13070__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_122_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08968_ _04312_ _01682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_87_Left_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07919_ _03160_ memory\[19\]\[11\] _03722_ _03724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08899_ _04231_ memory\[26\]\[23\] _04272_ _04276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10887__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10930_ _05383_ _00493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07752__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_158_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13125__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10861_ _05346_ _00461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12600_ _06322_ _06800_ _06461_ _06801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_112_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13580_ _05752_ _02967_ _05791_ _02968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_137_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13450__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10792_ _05043_ memory\[53\]\[18\] _05301_ _05310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12531_ _06446_ _06727_ _06730_ _06732_ _06733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__10367__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_96_Left_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15250_ _00209_ clknet_leaf_39_clk_i memory\[46\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13202__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12462_ _06322_ _06664_ _06461_ _06665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_10_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14201_ _01240_ clknet_leaf_108_clk_i memory\[19\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11413_ _03353_ memory\[62\]\[21\] _05638_ _05640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12582__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15181_ _00140_ clknet_leaf_386_clk_i memory\[44\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12556__A3 _06741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12393_ memory\[46\]\[12\] memory\[47\]\[12\] _06596_ _06597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07676__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14132_ _01171_ clknet_leaf_136_clk_i memory\[6\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10811__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11344_ _05603_ _00687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_61_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_84_clk_i clknet_5_17__leaf_clk_i clknet_leaf_84_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14063_ _01102_ clknet_leaf_203_clk_i memory\[10\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11275_ _05566_ _00655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_37_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13014_ _06720_ _02410_ _02411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XPHY_EDGE_ROW_148_Right_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_123_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10226_ _04623_ memory\[45\]\[23\] _04991_ _04995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11926__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_99_clk_i clknet_5_21__leaf_clk_i clknet_leaf_99_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_33_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10157_ _04958_ _00145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_33_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10088_ _04621_ memory\[43\]\[22\] _04919_ _04922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14965_ _02004_ clknet_leaf_73_clk_i memory\[37\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13916_ _00955_ clknet_leaf_285_clk_i memory\[8\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_22_clk_i clknet_5_5__leaf_clk_i clknet_leaf_22_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14896_ _01935_ clknet_leaf_76_clk_i memory\[35\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13847_ _00886_ clknet_leaf_111_clk_i memory\[13\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_18_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_18_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13778_ _00817_ clknet_leaf_120_clk_i memory\[14\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13441__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12875__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09131__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15517_ _00476_ clknet_leaf_344_clk_i memory\[55\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13161__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12729_ _06428_ _02122_ _02129_ _02130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_37_clk_i clknet_5_7__leaf_clk_i clknet_leaf_37_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_183_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11460__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_wire76_I _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15448_ _00407_ clknet_leaf_269_clk_i memory\[52\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_330 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11055__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09799__I1 _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15379_ _00338_ clknet_leaf_157_clk_i memory\[50\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07586__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09940_ _04843_ _00043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11507__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07385__I _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_115_Right_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09871_ _04608_ memory\[40\]\[16\] _04800_ _04807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09420__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_70_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08822_ _03196_ _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_174_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08210__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08753_ _04184_ _01595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07704_ _03144_ memory\[63\]\[6\] _03603_ _03610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10869__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08684_ _04147_ _01563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07734__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13680__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_71_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13107__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07635_ _03573_ _01088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_95_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13432__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07566_ _03536_ _01056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09041__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09305_ _04229_ memory\[32\]\[22\] _04488_ _04491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11294__I0 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_193_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_64_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07497_ _03499_ _01024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_153_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09976__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09236_ _04454_ _01808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08880__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09239__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_17_Right_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_170_3641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_90_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11046__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09167_ _04227_ memory\[30\]\[21\] _04416_ _04418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10915__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07496__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08118_ _03802_ memory\[15\]\[24\] _03841_ _03846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_133_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09098_ _04381_ _01743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08049_ _03806_ memory\[12\]\[26\] _03794_ _03807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07965__A3 _03123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13043__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11349__I1 _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11060_ _05452_ _00554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09411__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12171__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10011_ _04612_ memory\[42\]\[18\] _04872_ _04881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10650__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_26_Right_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_output57_I net57 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09216__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08120__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_188_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11545__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14750_ _01789_ clknet_leaf_412_clk_i memory\[31\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_4_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11962_ _06024_ _06167_ _06169_ _06171_ _06172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_157_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07725__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13701_ _03081_ _00768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10913_ memory\[55\]\[10\] _03155_ _05374_ _05375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14681_ _01720_ clknet_leaf_85_clk_i memory\[28\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11893_ memory\[38\]\[5\] memory\[39\]\[5\] _06039_ _06104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_39_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13632_ memory\[52\]\[31\] memory\[53\]\[31\] _05716_ _03019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13423__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10844_ _05026_ memory\[54\]\[10\] _05337_ _05338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_147_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_184_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13563_ _02950_ _02951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_67_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10775_ _05289_ _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_165_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08150__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_35_Right_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15302_ _00261_ clknet_leaf_294_clk_i memory\[48\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12514_ _06715_ _06716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09886__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12609__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13494_ _02367_ _02879_ _02881_ _02883_ _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_180_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15233_ _00192_ clknet_leaf_417_clk_i memory\[46\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12445_ _06647_ _06648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_151_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10825__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11737__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13201__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_508 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15164_ _00123_ clknet_leaf_421_clk_i memory\[44\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12376_ memory\[14\]\[12\] memory\[15\]\[12\] _06302_ _06580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_26_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_1_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14115_ _01154_ clknet_leaf_300_clk_i memory\[6\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11327_ _05594_ _00679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15095_ _00054_ clknet_leaf_10_clk_i memory\[41\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14046_ _01085_ clknet_leaf_309_clk_i memory\[10\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_52_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11258_ _05557_ _00647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_44_Right_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_52_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07169__A1 _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12162__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10560__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10209_ _04606_ memory\[45\]\[15\] _04980_ _04986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11189_ _03334_ memory\[5\]\[12\] _05518_ _05521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11455__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14948_ _01987_ clknet_leaf_431_clk_i memory\[37\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08965__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12487__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14879_ _01918_ clknet_leaf_424_clk_i memory\[35\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07192__I1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07420_ memory\[49\]\[2\] _03313_ _03455_ _03458_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_53_Right_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_67_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11276__I0 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07351_ _03419_ _00958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07282_ memory\[11\]\[3\] _03315_ _03379_ _03383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09021_ _04340_ _01707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11028__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10735__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13273__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11728__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09641__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_349_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_62_Right_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_141_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09923_ _04834_ _00035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09854_ _04591_ memory\[40\]\[8\] _04789_ _04798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10470__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08939__I _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08805_ _04219_ _01612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_146_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_146_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_401_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09785_ _04760_ _02051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06997_ _03203_ memory\[14\]\[25\] _03188_ _03204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08736_ _04174_ _01588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_107_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13653__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_1_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08667_ memory\[23\]\[25\] _03361_ _04132_ _04138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07183__I1 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_EDGE_ROW_71_Right_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_178_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07618_ _03563_ _01081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08598_ _03804_ memory\[22\]\[25\] _04095_ _04101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_37_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11267__I0 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07549_ _03526_ _01049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_48_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08132__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11511__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_147_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10560_ _05016_ memory\[50\]\[5\] _05181_ _05187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09880__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09219_ _04445_ _01800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12924__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10490__I1 memory\[4\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10491_ _05150_ _00287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_16_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11719__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12230_ _06155_ _06430_ _06433_ _06435_ _06436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__06922__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_32_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_32_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12145__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Right_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12161_ memory\[0\]\[9\] memory\[1\]\[9\] memory\[2\]\[9\] memory\[3\]\[9\] _06020_
+ _06090_ _06368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_31_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07954__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11112_ _03325_ memory\[58\]\[8\] _05471_ _05480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12092_ memory\[12\]\[8\] memory\[13\]\[8\] _06025_ _06300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_9_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_9_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11043_ _05443_ _00546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_73_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07946__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14802_ _01841_ clknet_leaf_76_clk_i memory\[32\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15782_ _00741_ clknet_leaf_254_clk_i net41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09699__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12994_ memory\[52\]\[21\] memory\[53\]\[21\] _06832_ _02391_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_93_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14733_ _01772_ clknet_leaf_127_clk_i memory\[30\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11945_ _05653_ _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_87_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08371__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07174__I1 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14664_ _01703_ clknet_leaf_181_clk_i memory\[28\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11876_ _06086_ _06087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_298_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13615_ _03002_ _03003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10827_ _05010_ memory\[54\]\[2\] _05326_ _05329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14595_ _01634_ clknet_leaf_409_clk_i memory\[26\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13546_ memory\[30\]\[29\] memory\[31\]\[29\] _05737_ _02935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10758_ _05292_ _00412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09871__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13477_ memory\[40\]\[28\] memory\[41\]\[28\] memory\[42\]\[28\] memory\[43\]\[28\]
+ _05692_ _05694_ _02867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_70_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10689_ _05008_ memory\[52\]\[1\] _05254_ _05256_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15216_ _00175_ clknet_leaf_17_clk_i memory\[45\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12428_ _06272_ _06626_ _06628_ _06630_ _06631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__09623__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_350_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15147_ _00106_ clknet_leaf_33_clk_i memory\[43\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_168_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12359_ memory\[52\]\[12\] memory\[53\]\[12\] _06143_ _06563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11894__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15078_ _00037_ clknet_leaf_29_clk_i memory\[41\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14029_ _01068_ clknet_leaf_170_clk_i memory\[0\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_06920_ _03145_ _00801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10290__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09570_ _04646_ _01950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08695__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13635__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_89 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08521_ _04060_ _01487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_141_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08452_ _03793_ memory\[20\]\[20\] _04023_ _04024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12010__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_65_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07403_ _03446_ _00983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08383_ _03964_ _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08114__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_84 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07334_ memory\[11\]\[28\] _03367_ _03401_ _03410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08665__I1 _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07265_ _03217_ _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_26_480 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09004_ _04331_ _01699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_84_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07196_ _03324_ _00898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_143_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11421__I0 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10264__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12680__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_130_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07774__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_148_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12126__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11296__S _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09906_ _04573_ memory\[41\]\[0\] _04825_ _04826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_6_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12677__A2 _06876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09837_ _04788_ _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11095__I _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07553__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09768_ memory\[3\]\[0\] _03110_ _04751_ _04752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_193_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_5_0__f_clk_i_I clknet_2_0_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08719_ _04165_ _01580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13524__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09699_ _04573_ memory\[38\]\[0\] _04714_ _04715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_14_Left_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_11730_ memory\[52\]\[3\] memory\[53\]\[3\] _05678_ _05943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06917__I net35 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10160__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_550 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11661_ _05874_ _05875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_83_328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08105__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13485__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13400_ _05777_ _02790_ _02791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_25_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_25_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10612_ _05068_ memory\[50\]\[30\] _05180_ _05214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14380_ _01419_ clknet_leaf_172_clk_i memory\[1\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11592_ _05660_ _05806_ _05665_ _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_25_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13331_ _05747_ _02718_ _02720_ _02722_ _02723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_106_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10375__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10543_ _05177_ _00312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13262_ memory\[4\]\[25\] memory\[5\]\[25\] _06845_ _02655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_49_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10474_ _05066_ memory\[48\]\[29\] _05131_ _05141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09605__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_23_Left_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12365__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15001_ _02040_ clknet_leaf_65_clk_i memory\[38\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11799__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13686__S _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12213_ memory\[52\]\[10\] memory\[53\]\[10\] _06143_ _06419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12590__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13193_ memory\[54\]\[24\] memory\[55\]\[24\] _02312_ _02587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_121_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_185_3938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07684__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07092__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12144_ memory\[62\]\[9\] memory\[63\]\[9\] _05868_ _06351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12075_ _06272_ _06275_ _06278_ _06282_ _06283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07919__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11026_ _03452_ _03490_ _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_99_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11934__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15834_ _00793_ clknet_leaf_386_clk_i memory\[9\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13617__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_32_Left_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_86_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12977_ _05759_ _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_15765_ _00724_ clknet_leaf_148_clk_i memory\[62\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08344__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12140__I1 net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_443_clk_i clknet_5_1__leaf_clk_i clknet_leaf_443_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_59_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11928_ _05669_ _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14716_ _01755_ clknet_leaf_391_clk_i memory\[30\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15696_ _00655_ clknet_leaf_162_clk_i memory\[60\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_86_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14647_ _01686_ clknet_leaf_79_clk_i memory\[27\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11859_ _06070_ _00735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12765__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07859__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14578_ _01617_ clknet_leaf_81_clk_i memory\[25\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09844__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_43_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_60_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13529_ memory\[36\]\[29\] memory\[37\]\[29\] _02338_ _02918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08272__A2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_41_Left_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07050_ _03228_ _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_126_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07594__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12108__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07952_ _03209_ memory\[19\]\[27\] _03733_ _03741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06903_ _03132_ memory\[14\]\[2\] _03126_ _03133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07883_ _03704_ _01205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08583__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_50_Left_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09622_ _04673_ _01975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_74_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10390__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09553_ _04635_ memory\[35\]\[29\] _04617_ _04636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_121_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08504_ _04051_ _01479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09484_ _03146_ _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_78_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08435_ _03777_ memory\[20\]\[12\] _04012_ _04015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_19_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_21_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08366_ _03978_ _01414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_22_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13387__A3 _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08638__I1 _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_189_4005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_50_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_878 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07317_ _03378_ _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_33_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08297_ _03775_ memory\[18\]\[11\] _03940_ _03942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_93 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09984__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07248_ memory\[39\]\[24\] _03359_ _03351_ _03360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_131_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12347__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__I1 memory\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07179_ _03131_ _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_44_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_246_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10190_ _04587_ memory\[45\]\[6\] _04969_ _04976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07009__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12900_ _06467_ _02291_ _02298_ _02299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__11953__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13880_ _00919_ clknet_leaf_19_clk_i memory\[39\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10381__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09224__S _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12831_ memory\[22\]\[18\] memory\[23\]\[18\] _06751_ _02231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08326__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11553__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15550_ _00509_ clknet_leaf_326_clk_i memory\[56\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10133__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12762_ _02162_ _00748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_189_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_16_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14501_ _01540_ clknet_leaf_362_clk_i memory\[23\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11713_ _05926_ _05927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_56_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_178_3797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15481_ _00440_ clknet_leaf_269_clk_i memory\[53\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12693_ memory\[16\]\[16\] memory\[17\]\[16\] memory\[18\]\[16\] memory\[19\]\[16\]
+ _06342_ _06485_ _02095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_14432_ _01471_ clknet_leaf_353_clk_i memory\[21\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_42_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11644_ _05788_ _05858_ _05792_ _05859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_42_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08629__I1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14363_ _01402_ clknet_leaf_27_clk_i memory\[18\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xinput16 data_i[18] net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_11575_ _03113_ _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_80_843 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput27 data_i[28] net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07301__I1 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput38 data_i[9] net38 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__09894__S _04811_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13314_ memory\[56\]\[26\] memory\[57\]\[26\] memory\[58\]\[26\] memory\[59\]\[26\]
+ _05711_ _02171_ _02706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_181_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10526_ _05050_ memory\[4\]\[21\] _05167_ _05169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14294_ _01333_ clknet_leaf_84_clk_i memory\[29\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12338__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13245_ _02638_ net56 _02382_ _02639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10833__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10457_ _05132_ _00271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_122_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12433__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07065__I0 _03178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08303__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13176_ _02371_ _02570_ _02373_ _02571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10388_ _05047_ memory\[47\]\[20\] _05095_ _05096_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12127_ memory\[24\]\[8\] memory\[25\]\[8\] memory\[26\]\[8\] memory\[27\]\[8\] _05778_
+ _05922_ _06335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_97_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12058_ _05794_ _06266_ _06267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12510__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11009_ _05425_ _00530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15817_ _00776_ clknet_leaf_211_clk_i memory\[9\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13164__B _02556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_382_clk_i clknet_5_7__leaf_clk_i clknet_leaf_382_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_137_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08973__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10124__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15748_ _00707_ clknet_leaf_304_clk_i memory\[62\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10675__I1 _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12495__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15679_ _00638_ clknet_leaf_334_clk_i memory\[60\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07540__I1 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08220_ _03766_ memory\[17\]\[7\] _03893_ _03901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_397_clk_i clknet_5_3__leaf_clk_i clknet_leaf_397_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_195_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08772__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13369__A3 _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12577__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08151_ _03864_ _01313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_99_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07102_ _03269_ _00859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_320_clk_i clknet_5_11__leaf_clk_i clknet_leaf_320_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_71_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08082_ _03766_ memory\[15\]\[7\] _03819_ _03827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07033_ _03231_ _00828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10743__S _05276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09309__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_987 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_335_clk_i clknet_5_10__leaf_clk_i clknet_leaf_335_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08984_ _04320_ _01690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07935_ _03184_ memory\[19\]\[19\] _03722_ _03732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08556__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11574__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07866_ _03695_ _01197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09605_ _04616_ memory\[36\]\[20\] _04664_ _04665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input19_I data_i[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07797_ _03181_ memory\[6\]\[18\] _03650_ _03659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_27_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09536_ _04624_ _01938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_149_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire73 _03227_ net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09467_ _04577_ memory\[35\]\[1\] _04575_ _04578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08418_ _03760_ memory\[20\]\[4\] _04001_ _04006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08682__I _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09398_ _04540_ _01884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08349_ _03969_ _01406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_129_Right_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_11_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11360_ _05611_ _00695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10311_ _03190_ _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_11291_ _05574_ _00663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12415__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_397_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13030_ _02209_ _02422_ _02424_ _02426_ _02427_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__06930__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10242_ _04639_ memory\[45\]\[31\] _04968_ _05003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08795__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12740__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10173_ _04966_ _00153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14981_ _02020_ clknet_leaf_404_clk_i memory\[38\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13932_ _00971_ clknet_leaf_213_clk_i memory\[8\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10354__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13863_ _00902_ clknet_leaf_259_clk_i memory\[39\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15602_ _00561_ clknet_leaf_164_clk_i memory\[57\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12814_ memory\[46\]\[18\] memory\[47\]\[18\] _06596_ _02214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10106__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13794_ _00833_ clknet_leaf_340_clk_i memory\[16\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_1065 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_106_Left_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_69_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12745_ memory\[28\]\[17\] memory\[29\]\[17\] _06604_ _02146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15533_ _00492_ clknet_leaf_241_clk_i memory\[55\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_127_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15464_ _00423_ clknet_leaf_296_clk_i memory\[53\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12676_ memory\[40\]\[16\] memory\[41\]\[16\] memory\[42\]\[16\] memory\[43\]\[16\]
+ _06875_ _06326_ _06876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XFILLER_0_127_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12328__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14415_ _01454_ clknet_leaf_188_clk_i memory\[20\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11627_ _05841_ _05842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_182_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15395_ _00354_ clknet_leaf_334_clk_i memory\[51\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_13_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13220__A2 _02609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14346_ _01385_ clknet_leaf_207_clk_i memory\[18\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11558_ memory\[30\]\[0\] memory\[31\]\[0\] _05773_ _05774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10509_ _05033_ memory\[4\]\[13\] _05156_ _05160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14277_ _01316_ clknet_leaf_360_clk_i memory\[29\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11489_ _05659_ _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__13603__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09129__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07038__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_94_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13228_ _02336_ _02614_ _02621_ _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_21_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08786__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_55_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_55_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13159_ _02553_ _02554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07872__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_72_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08538__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11394__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07720_ _03618_ _01128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11917__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11298__A1 _03266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07651_ _03166_ memory\[10\]\[13\] _03578_ _03582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10896__I1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09799__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07582_ _03166_ memory\[0\]\[13\] _03541_ _03545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_125_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12798__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09321_ _04245_ memory\[32\]\[30\] _04465_ _04499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10648__I1 _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08710__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07513__I1 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09252_ _04462_ _01816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08208__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08203_ _03891_ _01338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09183_ _04243_ memory\[30\]\[29\] _04416_ _04426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12953__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08134_ _03113_ _03224_ _03854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_116_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_940 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_151_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08065_ _03817_ _01274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_109_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_112_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09039__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07016_ _03217_ _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__13069__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_274_clk_i clknet_5_13__leaf_clk_i clknet_leaf_274_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_112_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_773 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13070__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11368__I _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08878__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08967_ _04231_ memory\[27\]\[23\] _04308_ _04312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_289_clk_i clknet_5_15__leaf_clk_i clknet_leaf_289_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07918_ _03723_ _01221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10336__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08898_ _04275_ _01649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07849_ _03156_ memory\[7\]\[10\] _03686_ _03687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_3_clk_i clknet_5_4__leaf_clk_i clknet_leaf_3_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_212_clk_i clknet_5_30__leaf_clk_i clknet_leaf_212_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10860_ _05043_ memory\[54\]\[18\] _05337_ _05346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12789__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_184_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09519_ _04612_ memory\[35\]\[18\] _04596_ _04613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13532__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10791_ _05309_ _00428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10648__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08701__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07504__I1 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13024__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12530_ _06453_ _06731_ _06732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_109_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06925__I net37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08118__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_35_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_227_clk_i clknet_5_26__leaf_clk_i clknet_leaf_227_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_53_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12461_ memory\[46\]\[13\] memory\[47\]\[13\] _06596_ _06664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12863__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14200_ _01239_ clknet_leaf_110_clk_i memory\[19\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_152_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11412_ _05639_ _00719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15180_ _00139_ clknet_leaf_37_clk_i memory\[44\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12392_ _05701_ _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12556__A4 _06757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14131_ _01170_ clknet_leaf_119_clk_i memory\[6\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11343_ memory\[61\]\[20\] _03186_ _05602_ _05603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10383__S _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14062_ _01101_ clknet_leaf_204_clk_i memory\[10\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11274_ _03350_ memory\[60\]\[20\] _05565_ _05566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13013_ memory\[8\]\[21\] memory\[9\]\[21\] memory\[10\]\[21\] memory\[11\]\[21\]
+ _06582_ _06721_ _02410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__13694__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12713__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10225_ _04994_ _00177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_143_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10575__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07692__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10156_ _04621_ memory\[44\]\[22\] _04955_ _04958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_33_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12611__B _06809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08587__I _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10087_ _04921_ _00112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10327__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14964_ _02003_ clknet_leaf_12_clk_i memory\[37\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09193__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13915_ _00954_ clknet_leaf_387_clk_i memory\[11\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14895_ _01934_ clknet_leaf_63_clk_i memory\[35\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08940__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13846_ _00885_ clknet_leaf_110_clk_i memory\[13\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_18_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13777_ _00816_ clknet_leaf_113_clk_i memory\[14\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10558__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10989_ _05035_ memory\[56\]\[14\] _05410_ _05415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_29_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12875__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15516_ _00475_ clknet_leaf_332_clk_i memory\[55\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12728_ _06713_ _02124_ _02126_ _02128_ _02129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_17_309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_618 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09211__I _04429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_68_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12659_ memory\[8\]\[16\] memory\[9\]\[16\] memory\[10\]\[16\] memory\[11\]\[16\]
+ _06582_ _06721_ _06859_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_15447_ _00406_ clknet_leaf_268_clk_i memory\[52\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_167_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07867__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_96_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15378_ _00337_ clknet_leaf_157_clk_i memory\[50\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_111_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14329_ _01368_ clknet_leaf_106_clk_i memory\[17\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_57_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10293__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_74_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13752__I0 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09870_ _04806_ _00010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10566__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_7__f_clk_i clknet_2_0_0_clk_i clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08821_ _04230_ _01617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13617__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08752_ _04181_ memory\[25\]\[0\] _04183_ _04184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10318__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08136__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07703_ _03609_ _01120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07107__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12563__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08683_ _03746_ memory\[24\]\[0\] _04146_ _04147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08931__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07634_ _03141_ memory\[10\]\[5\] _03567_ _03573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_345_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07565_ _03141_ memory\[0\]\[5\] _03530_ _03536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10468__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_49_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_192_4067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09304_ _04490_ _01840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07496_ memory\[59\]\[5\] _03319_ _03493_ _03499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_153_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_153_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09235_ _04227_ memory\[31\]\[21\] _04452_ _04454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_746 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12683__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10267__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13196__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09166_ _04417_ _01775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08960__I _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_160_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08117_ _03845_ _01298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_131_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09097_ _04224_ memory\[2\]\[20\] _04380_ _04381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09992__S _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07670__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08048_ _03205_ _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_43_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_31_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13043__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10931__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10010_ _04880_ _00076_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09999_ _04600_ memory\[42\]\[12\] _04872_ _04875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13019__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10309__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07017__S _03125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_4_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11961_ _06031_ _06170_ _06171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12858__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_151_clk_i clknet_5_19__leaf_clk_i clknet_leaf_151_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_4_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11762__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_1249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13700_ _03319_ memory\[9\]\[5\] _03075_ _03081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10912_ _05362_ _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14680_ _01719_ clknet_leaf_85_clk_i memory\[28\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11682__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11892_ _06102_ _06103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_86_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13631_ _05700_ _03013_ _03015_ _03017_ _03018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10843_ _05325_ _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11561__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_166_clk_i clknet_5_25__leaf_clk_i clknet_leaf_166_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13562_ memory\[60\]\[30\] memory\[61\]\[30\] _05702_ _02950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10774_ _05300_ _00420_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_54_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_181_Right_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12513_ memory\[12\]\[14\] memory\[13\]\[14\] _06714_ _06715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15301_ _00260_ clknet_leaf_317_clk_i memory\[48\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10177__I _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13493_ _02375_ _02882_ _02883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12609__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_168_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13187__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12444_ memory\[12\]\[13\] memory\[13\]\[13\] _06025_ _06647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15232_ _00191_ clknet_leaf_417_clk_i memory\[46\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08989__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15163_ _00122_ clknet_leaf_441_clk_i memory\[43\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12392__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12375_ _06578_ _06579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_1_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11002__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14114_ _01153_ clknet_leaf_300_clk_i memory\[6\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07661__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11326_ memory\[61\]\[12\] _03162_ _05591_ _05594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15094_ _00053_ clknet_leaf_6_clk_i memory\[41\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_91_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11937__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13734__I0 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14045_ _01084_ clknet_leaf_288_clk_i memory\[10\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_104_clk_i clknet_5_21__leaf_clk_i clknet_leaf_104_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10841__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11257_ _03334_ memory\[60\]\[12\] _05554_ _05557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_294_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_52_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07169__A2 _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09407__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12162__A2 _06368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10208_ _04985_ _00169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08311__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11188_ _05520_ _00614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_59_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10139_ _04604_ memory\[44\]\[14\] _04944_ _04949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_94_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_119_clk_i clknet_5_23__leaf_clk_i clknet_leaf_119_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12768__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14947_ _01986_ clknet_leaf_432_clk_i memory\[37\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08913__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_1304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11673__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14878_ _01917_ clknet_leaf_424_clk_i memory\[35\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10720__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13829_ _00868_ clknet_leaf_288_clk_i memory\[13\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11471__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_147_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07350_ _03135_ memory\[8\]\[3\] _03415_ _03419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08981__S _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_31_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13599__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07281_ _03382_ _00925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_73_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13178__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09020_ _04216_ memory\[28\]\[16\] _04333_ _04340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07597__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_122_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_72_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_470 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13273__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12008__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13725__I0 _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09922_ _04591_ memory\[41\]\[8\] _04825_ _04834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10751__S _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07404__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09853_ _04797_ _00002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08804_ _04218_ memory\[25\]\[17\] _04204_ _04219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_146_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09784_ memory\[3\]\[8\] _03149_ _04751_ _04760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_146_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06996_ _03202_ _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__12536__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08020__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08735_ _03804_ memory\[24\]\[25\] _04168_ _04174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_107_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_107_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_1_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08666_ _04137_ _01555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_124_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_83_clk_i clknet_5_20__leaf_clk_i clknet_leaf_83_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_178_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07617_ _03218_ memory\[0\]\[30\] _03529_ _03563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08597_ _04100_ _01523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_193_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07548_ memory\[59\]\[30\] _03371_ _03492_ _03526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11511__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_162_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_884 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07479_ _03488_ _01017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_640 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_98_clk_i clknet_5_21__leaf_clk_i clknet_leaf_98_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13169__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09218_ _04210_ memory\[31\]\[13\] _04441_ _04445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10490_ _05014_ memory\[4\]\[4\] _05145_ _05150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_45_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12916__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09149_ _04408_ _01767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10778__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_21_clk_i clknet_5_5__leaf_clk_i clknet_leaf_21_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12160_ _06159_ _06366_ _06018_ _06367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_124_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11111_ _05479_ _00578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12940__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12091_ _06155_ _06294_ _06296_ _06298_ _06299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_102_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10661__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_9_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11042_ _05020_ memory\[57\]\[7\] _05435_ _05443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_16_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13257__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11556__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_183_3888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_36_clk_i clknet_5_7__leaf_clk_i clknet_leaf_36_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_183_3899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09148__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14801_ _01840_ clknet_leaf_61_clk_i memory\[32\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15781_ _00740_ clknet_leaf_338_clk_i net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12993_ _02163_ _02385_ _02387_ _02389_ _02390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_118_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14732_ _01771_ clknet_leaf_127_clk_i memory\[30\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_99_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11944_ _05651_ _06141_ _06153_ _06154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_98_164 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_118_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14663_ _01702_ clknet_leaf_177_clk_i memory\[28\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11875_ memory\[4\]\[5\] memory\[5\]\[5\] _05702_ _06086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10826_ _05328_ _00444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13614_ memory\[20\]\[30\] memory\[21\]\[30\] _05749_ _03002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14594_ _01633_ clknet_leaf_409_clk_i memory\[26\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_32_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_82_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13545_ _02933_ _02934_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10757_ _05008_ memory\[53\]\[1\] _05290_ _05292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12080__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07882__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13476_ _05682_ _02865_ _02352_ _02866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10688_ _05255_ _00379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12336__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15215_ _00174_ clknet_leaf_34_clk_i memory\[45\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12427_ _06279_ _06629_ _06630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_124_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10769__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13580__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07634__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15146_ _00105_ clknet_leaf_21_clk_i memory\[43\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12358_ _06272_ _06556_ _06559_ _06561_ _06562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_10_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11309_ memory\[61\]\[4\] _03137_ _05580_ _05585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15077_ _00036_ clknet_leaf_431_clk_i memory\[41\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10571__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_25__f_clk_i clknet_2_3_0_clk_i clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12289_ _06493_ _06494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_77_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09387__I0 _04243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14028_ _01067_ clknet_leaf_171_clk_i memory\[0\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09137__S _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11466__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11894__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07880__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09139__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08520_ _03793_ memory\[21\]\[20\] _04059_ _04060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_5_30__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11646__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08775__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08451_ _04000_ _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07402_ _03212_ memory\[8\]\[28\] _03437_ _03446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08382_ _03986_ _01422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_45_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09600__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09311__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07333_ _03409_ _00950_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07264_ _03370_ _00920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08216__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09003_ _04199_ memory\[28\]\[8\] _04322_ _04331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12246__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_604 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12961__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07195_ memory\[39\]\[7\] _03323_ _03309_ _03324_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_13_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_83_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09047__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13323__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09905_ _04824_ _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_165_3552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11185__I0 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10280__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09836_ net73 _04787_ _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08886__S _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08750__A1 net74 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_77_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09767_ _04750_ _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_06979_ net20 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_154_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08718_ _03787_ memory\[24\]\[17\] _04157_ _04165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11637__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09698_ _04713_ _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_55_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09550__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08649_ _04128_ _01547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_242_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_84_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_138_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11660_ memory\[52\]\[2\] memory\[53\]\[2\] _05678_ _05874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_154_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09510__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13485__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_25_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10611_ _05213_ _00344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_25_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11496__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11591_ memory\[62\]\[1\] memory\[63\]\[1\] _05662_ _05806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10656__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10999__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13032__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13330_ _05759_ _02721_ _02722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_14_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_106_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06933__I net8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10542_ _05066_ memory\[4\]\[29\] _05167_ _05177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08126__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07030__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_464 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13261_ _02302_ _02646_ _02653_ _02654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_17_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10455__I _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10473_ _05140_ _00279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12871__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15000_ _02039_ clknet_leaf_19_clk_i memory\[38\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12212_ _06272_ _06413_ _06415_ _06417_ _06418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_121_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11799__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13192_ _02585_ _02586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_185_3928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11487__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12143_ _06349_ _06350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_23_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09369__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12074_ _06279_ _06281_ _06282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11176__I0 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11025_ _05433_ _00538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15833_ _00792_ clknet_leaf_132_clk_i memory\[9\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_86_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15764_ _00723_ clknet_leaf_147_clk_i memory\[62\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12976_ _02371_ _02372_ _02373_ _02374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_47_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09541__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14715_ _01754_ clknet_leaf_28_clk_i memory\[2\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11927_ _05660_ _06136_ _06001_ _06137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15695_ _00654_ clknet_leaf_255_clk_i memory\[60\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11950__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14646_ _01685_ clknet_leaf_82_clk_i memory\[27\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11858_ _06069_ net66 _05802_ _06070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_74_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07004__I _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_83_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09420__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10566__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10809_ _05060_ memory\[53\]\[26\] _05312_ _05319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14577_ _01616_ clknet_leaf_93_clk_i memory\[25\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11100__I0 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11789_ _05664_ _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_60_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07855__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13528_ _02319_ _02909_ _02916_ _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_27_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11800__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13459_ _02848_ _02849_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_141_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_444_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07607__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08280__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15129_ _00088_ clknet_leaf_7_clk_i memory\[42\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13305__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_189_Left_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07951_ _03740_ _01237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_191_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06902_ _03131_ _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_07882_ _03206_ memory\[7\]\[26\] _03697_ _03704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_143_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_09621_ _04633_ memory\[36\]\[28\] _04664_ _04673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_160_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09552_ _03214_ _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XTAP_TAPCELL_ROW_121_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08503_ _03777_ memory\[21\]\[12\] _04048_ _04051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07115__S _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09532__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09483_ _04588_ _01921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11860__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08434_ _04014_ _01446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08099__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12044__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08365_ _03775_ memory\[1\]\[11\] _03976_ _03978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10476__S _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07316_ _03400_ _00942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_189_4017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_149_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07846__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08296_ _03941_ _01381_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_119_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07247_ _03199_ _03359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_119_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12691__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12347__A2 _06544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07785__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07178_ _03312_ _00892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11100__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11158__I0 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_180_3836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_180_3847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09819_ _04778_ _02067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11953__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13155__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12830_ _02229_ _02230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12283__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12761_ _02161_ net48 _06491_ _02162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_393_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11770__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14500_ _01539_ clknet_leaf_362_clk_i memory\[23\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11712_ memory\[20\]\[2\] memory\[21\]\[2\] _05785_ _05926_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_178_3798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12692_ _06480_ _02093_ _06482_ _02094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15480_ _00439_ clknet_leaf_380_clk_i memory\[53\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14431_ _01470_ clknet_leaf_353_clk_i memory\[21\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11643_ memory\[22\]\[1\] memory\[23\]\[1\] _05789_ _05858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_42_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09826__I1 _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07759__I _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11574_ memory\[22\]\[0\] memory\[23\]\[0\] _05789_ _05790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14362_ _01401_ clknet_leaf_26_clk_i memory\[18\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput17 data_i[19] net17 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
Xinput28 data_i[29] net28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_10525_ _05168_ _00303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13313_ _02167_ _02704_ _05756_ _02705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
Xinput39 we_i net39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_14293_ _01332_ clknet_leaf_83_clk_i memory\[29\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_162_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13244_ _02592_ _02607_ _02622_ _02637_ _02638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_10456_ _05047_ memory\[48\]\[20\] _05131_ _05132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_161_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13175_ memory\[22\]\[23\] memory\[23\]\[23\] _06751_ _02570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08262__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10387_ _05072_ _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11010__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12126_ _05918_ _06333_ _06195_ _06334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_97_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12057_ memory\[16\]\[7\] memory\[17\]\[7\] memory\[18\]\[7\] memory\[19\]\[7\] _05795_
+ _05796_ _06266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12510__A2 _06705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11008_ _05054_ memory\[56\]\[23\] _05421_ _05425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15816_ _00775_ clknet_leaf_210_clk_i memory\[9\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15747_ _00706_ clknet_leaf_304_clk_i memory\[62\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_88_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12959_ _02336_ _02348_ _02356_ _02357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_15678_ _00637_ clknet_leaf_327_clk_i memory\[60\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09150__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_138_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12026__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14629_ _01668_ clknet_leaf_408_clk_i memory\[27\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10296__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08150_ _03764_ memory\[29\]\[6\] _03857_ _03864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07828__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07101_ _03111_ memory\[13\]\[0\] _03268_ _03269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_99_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08081_ _03826_ _01281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_153_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13526__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07032_ _03129_ memory\[16\]\[1\] _03229_ _03231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_141_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12016__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_114_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10060__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08983_ _04247_ memory\[27\]\[31\] _04285_ _04320_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_110_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07934_ _03731_ _01229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09753__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07865_ _03181_ memory\[7\]\[18\] _03686_ _03695_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11654__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09604_ _04641_ _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_190_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07796_ _03658_ _01164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12265__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_27_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09535_ _04623_ memory\[35\]\[23\] _04617_ _04624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_167_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09466_ _03128_ _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_4_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_94_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08417_ _04005_ _01438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09397_ _04185_ memory\[34\]\[1\] _04538_ _04540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09995__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08348_ _03758_ memory\[1\]\[3\] _03965_ _03969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08492__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08279_ _03932_ _01373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10934__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11871__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13310__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13517__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10310_ _05049_ _00207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_116_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11290_ _03367_ memory\[60\]\[28\] _05565_ _05574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08404__S _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11379__I0 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10241_ _05002_ _00185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11623__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_442_clk_i clknet_5_1__leaf_clk_i clknet_leaf_442_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09992__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12740__A2 _02140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10172_ _04637_ memory\[44\]\[30\] _04932_ _04966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14980_ _02019_ clknet_leaf_401_clk_i memory\[38\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09235__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13931_ _00970_ clknet_leaf_210_clk_i memory\[8\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13265__B _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13862_ _00901_ clknet_leaf_272_clk_i memory\[39\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15601_ _00560_ clknet_leaf_165_clk_i memory\[57\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12256__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12813_ _05681_ _02213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_13793_ _00832_ clknet_leaf_343_clk_i memory\[16\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09121__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15532_ _00491_ clknet_leaf_241_clk_i memory\[55\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12744_ _06445_ _02137_ _02144_ _02145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_15463_ _00422_ clknet_leaf_295_clk_i memory\[53\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12675_ _05691_ _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_155_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14414_ _01453_ clknet_leaf_190_clk_i memory\[20\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11626_ memory\[44\]\[1\] memory\[45\]\[1\] _05749_ _05841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_25_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15394_ _00353_ clknet_leaf_313_clk_i memory\[51\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_142_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14345_ _01384_ clknet_leaf_206_clk_i memory\[18\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07286__I1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11557_ _05683_ _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10844__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10290__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_52_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10508_ _05159_ _00295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14276_ _01315_ clknet_leaf_377_clk_i memory\[29\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11488_ _05703_ _05704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_123_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13603__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08235__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13227_ _02209_ _02616_ _02618_ _02620_ _02621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_94_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10439_ _05031_ memory\[48\]\[12\] _05120_ _05123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10042__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_55_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13158_ memory\[44\]\[23\] memory\[45\]\[23\] _02210_ _02553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_55_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11675__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_10 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12109_ _05732_ _06311_ _06313_ _06316_ _06317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_13089_ memory\[44\]\[22\] memory\[45\]\[22\] _02210_ _02485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_72_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_64_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11917__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11298__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_109_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11474__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07650_ _03581_ _01095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07581_ _03544_ _01063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09879__I _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09320_ _04498_ _01848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12798__A2 _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09251_ _04243_ memory\[31\]\[29\] _04452_ _04462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_289_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_138_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_28_351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08202_ _03816_ memory\[29\]\[31\] _03856_ _03891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09182_ _04425_ _01783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08133_ _03853_ _01306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_79_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_16_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_79_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08474__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11853__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13130__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10281__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08064_ _03816_ memory\[12\]\[31\] _03751_ _03817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08224__S _03893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_341_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07015_ net30 _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_109_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_112_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09974__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08023__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08966_ _04311_ _01681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_input31_I data_i[31] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09055__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09726__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07917_ _03156_ memory\[19\]\[10\] _03722_ _03723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13085__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08897_ _04229_ memory\[26\]\[22\] _04272_ _04275_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07201__I1 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07848_ _03674_ _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_162_Right_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12238__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10929__S _05374_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06960__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07779_ _03649_ _01156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09518_ _03180_ _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_39_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10790_ _05041_ memory\[53\]\[17\] _05301_ _05309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_175_3735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07303__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10728__I _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09449_ _04237_ memory\[34\]\[26\] _04560_ _04567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_192_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_163_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12460_ _06662_ _06663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_163_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_10_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11411_ _03350_ memory\[62\]\[20\] _05638_ _05639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12410__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12391_ _06594_ _06595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12943__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14130_ _01169_ clknet_leaf_119_clk_i memory\[6\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_22_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11342_ _05579_ _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_61_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_381_clk_i clknet_5_7__leaf_clk_i clknet_leaf_381_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11559__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14061_ _01100_ clknet_leaf_204_clk_i memory\[10\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11273_ _05542_ _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_123_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08917__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10024__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13012_ _06717_ _02408_ _02195_ _02409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10224_ _04621_ memory\[45\]\[22\] _04991_ _04994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10155_ _04957_ _00144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_396_clk_i clknet_5_3__leaf_clk_i clknet_leaf_396_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09717__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12477__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10086_ _04619_ memory\[43\]\[21\] _04919_ _04921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14963_ _02002_ clknet_leaf_73_clk_i memory\[37\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_50_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13914_ _00953_ clknet_leaf_386_clk_i memory\[11\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14894_ _01933_ clknet_leaf_64_clk_i memory\[35\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12229__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_13845_ _00884_ clknet_leaf_112_clk_i memory\[13\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10839__S _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_18_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08309__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13776_ _00815_ clknet_leaf_121_clk_i memory\[14\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10988_ _05414_ _00520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_290_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15515_ _00474_ clknet_leaf_376_clk_i memory\[54\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12727_ _06720_ _02127_ _02128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
Xclkbuf_leaf_334_clk_i clknet_5_10__leaf_clk_i clknet_leaf_334_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_127_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15446_ _00405_ clknet_leaf_267_clk_i memory\[52\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12658_ _06717_ _06857_ _06304_ _06858_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_44_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07012__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08456__I0 _03798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_866 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11609_ _05710_ _05823_ _05824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_167_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15377_ _00336_ clknet_leaf_156_clk_i memory\[50\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12589_ _06428_ _06782_ _06789_ _06790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_68_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14328_ _01367_ clknet_leaf_107_clk_i memory\[17\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_349_clk_i clknet_5_8__leaf_clk_i clknet_leaf_349_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_57_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08208__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14259_ _01298_ clknet_leaf_116_clk_i memory\[15\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_150_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08979__S _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09956__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_08820_ _04229_ memory\[25\]\[22\] _04225_ _04230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08778__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12012__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08751_ _04182_ _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07702_ _03141_ memory\[63\]\[5\] _03603_ _03609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12563__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08682_ _04145_ _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_109_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07633_ _03572_ _01087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10749__S _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11932__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07564_ _03535_ _01055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_193_716 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_192_4057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13432__A3 _02822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_4068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09303_ _04227_ memory\[32\]\[21\] _04488_ _04490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08695__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07495_ _03498_ _01023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07498__I1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09234_ _04453_ _01807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_153_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_3_Right_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_111_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_125_Left_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_56_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1085 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08447__I0 _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09165_ _04224_ memory\[30\]\[20\] _04416_ _04417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12763__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10484__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08116_ _03800_ memory\[15\]\[23\] _03841_ _03845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_9_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_131_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09096_ _04357_ _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_131_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08047_ _03805_ _01268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10283__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07793__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07422__I1 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12171__A3 _06377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_134_Left_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09998_ _04874_ _00070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08949_ _04302_ _01673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_129_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11960_ memory\[8\]\[6\] memory\[9\]\[6\] memory\[10\]\[6\] memory\[11\]\[6\] _05893_
+ _06032_ _06170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_192_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_4_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_4_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_93_1254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09513__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10911_ _05373_ _00484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12938__I _03304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11891_ memory\[36\]\[5\] memory\[37\]\[5\] _05733_ _06102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13630_ _05710_ _03016_ _03017_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__13503__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_15_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10842_ _05336_ _00452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13561_ _02949_ _00760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10773_ _05024_ memory\[53\]\[9\] _05290_ _05300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_143_Left_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA_clkbuf_leaf_12_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15300_ _00259_ clknet_leaf_317_clk_i memory\[48\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_66_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12512_ _05677_ _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_180_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13492_ memory\[16\]\[28\] memory\[17\]\[28\] memory\[18\]\[28\] memory\[19\]\[28\]
+ _05761_ _02376_ _02882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_137_676 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15231_ _00190_ clknet_leaf_417_clk_i memory\[46\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_180_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12443_ _06155_ _06641_ _06643_ _06645_ _06646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_48_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10394__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15162_ _00121_ clknet_leaf_441_clk_i memory\[43\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12374_ memory\[12\]\[12\] memory\[13\]\[12\] _06025_ _06578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_105_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12490__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14113_ _01152_ clknet_leaf_300_clk_i memory\[6\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11325_ _05593_ _00678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_160_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15093_ _00052_ clknet_leaf_10_clk_i memory\[41\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_532 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_91_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14044_ _01083_ clknet_leaf_285_clk_i memory\[10\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11256_ _05556_ _00646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_237_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_152_Left_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_24_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_52_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10207_ _04604_ memory\[45\]\[14\] _04980_ _04985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08610__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11187_ _03332_ memory\[5\]\[11\] _05518_ _05520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10138_ _04948_ _00136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_20__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14946_ _01985_ clknet_leaf_433_clk_i memory\[37\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10069_ _04602_ memory\[43\]\[13\] _04908_ _04912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_89_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07007__I net27 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12870__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14877_ _01916_ clknet_leaf_429_clk_i memory\[35\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11673__A2 _05886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13828_ _00867_ clknet_leaf_276_clk_i memory\[13\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_273_clk_i clknet_5_13__leaf_clk_i clknet_leaf_273_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_161_Left_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_58_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12784__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13759_ _00798_ clknet_leaf_281_clk_i memory\[14\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07878__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10484__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07280_ memory\[11\]\[2\] _03313_ _03379_ _03382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_26_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15429_ _00388_ clknet_leaf_318_clk_i memory\[52\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_14_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_288_clk_i clknet_5_15__leaf_clk_i clknet_leaf_288_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_170_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10236__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07101__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_clk_i clknet_5_4__leaf_clk_i clknet_leaf_2_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_170_Left_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_211_clk_i clknet_5_27__leaf_clk_i clknet_leaf_211_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_145_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09929__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09921_ _04833_ _00034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13628__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09852_ _04589_ memory\[40\]\[7\] _04789_ _04797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08803_ _03177_ _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_146_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09783_ _04759_ _02050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_146_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_226_clk_i clknet_5_26__leaf_clk_i clknet_leaf_226_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_06995_ net24 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08734_ _04173_ _01587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12536__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_107_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09333__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_439_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08665_ memory\[23\]\[24\] _03359_ _04132_ _04137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12861__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06915__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07616_ _03562_ _01080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_89_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08596_ _03802_ memory\[22\]\[24\] _04095_ _04100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_48_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07547_ _03525_ _01048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_193_546 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_119_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_48_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_186_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07478_ memory\[49\]\[30\] _03371_ _03454_ _03488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09217_ _04444_ _01799_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_17_652 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09148_ _04208_ memory\[30\]\[12\] _04405_ _04408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09079_ _04371_ _01734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10942__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11110_ _03323_ memory\[58\]\[7\] _05471_ _05479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_187_3970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12090_ _06162_ _06297_ _06298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_31_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08412__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11041_ _05442_ _00545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_9_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_183_3889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10950__I1 _03211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_14800_ _01839_ clknet_leaf_77_clk_i memory\[32\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_157_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15780_ _00739_ clknet_leaf_338_clk_i net70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07159__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12992_ _02170_ _02388_ _02389_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_99_644 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09243__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14731_ _01770_ clknet_leaf_130_clk_i memory\[30\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_19_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11943_ _06142_ _06145_ _06148_ _06152_ _06153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_87_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11572__I _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14662_ _01701_ clknet_leaf_177_clk_i memory\[28\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11874_ _05651_ _06077_ _06084_ _06085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_184_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13613_ _02494_ _02996_ _02998_ _03000_ _03001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_71_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10825_ _05008_ memory\[54\]\[1\] _05326_ _05328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_1322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__12604__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14593_ _01632_ clknet_leaf_416_clk_i memory\[26\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_39_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07698__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10466__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13544_ memory\[28\]\[29\] memory\[29\]\[29\] _02495_ _02933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_45_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10756_ _05291_ _00411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_94_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_484 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13475_ memory\[46\]\[28\] memory\[47\]\[28\] _02487_ _02865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_180_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10687_ _05004_ memory\[52\]\[0\] _05254_ _05255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_164_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15214_ _00173_ clknet_leaf_34_clk_i memory\[45\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_35_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12426_ memory\[56\]\[13\] memory\[57\]\[13\] memory\[58\]\[13\] memory\[59\]\[13\]
+ _06138_ _06280_ _06629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09084__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_785 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15145_ _00104_ clknet_leaf_25_clk_i memory\[43\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10852__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12357_ _06279_ _06560_ _06561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_11_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09418__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11308_ _05584_ _00670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_388_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08322__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15076_ _00035_ clknet_leaf_442_clk_i memory\[41\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12288_ memory\[60\]\[11\] memory\[61\]\[11\] _06273_ _06493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14027_ _01066_ clknet_leaf_218_clk_i memory\[0\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11239_ _05547_ _00638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07398__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13096__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_69_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_136_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_440_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12578__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14929_ _01968_ clknet_leaf_18_clk_i memory\[36\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10299__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08450_ _04022_ _01454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_373 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07401_ _03445_ _00982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08381_ _03791_ memory\[1\]\[19\] _03976_ _03986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_102_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_46_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07332_ memory\[11\]\[27\] _03365_ _03401_ _03409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13403__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08791__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_85_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_128_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07263_ memory\[39\]\[29\] _03369_ _03351_ _03370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09002_ _04330_ _01698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10209__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07194_ _03146_ _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_60_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07200__I _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_150_clk_i clknet_5_19__leaf_clk_i clknet_leaf_150_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11858__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11582__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13358__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_148_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_148_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09904_ net74 _04787_ _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_10_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_6_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_165_clk_i clknet_5_28__leaf_clk_i clknet_leaf_165_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09835_ _04786_ _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__12689__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09766_ _04749_ _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_06978_ _03189_ _00815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_20_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09063__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08717_ _04164_ _01579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13093__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12488__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09697_ _03124_ _03305_ _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_83_91 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08648_ memory\[23\]\[16\] _03342_ _04121_ _04128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07561__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08579_ _03785_ memory\[22\]\[16\] _04084_ _04091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_103_clk_i clknet_5_21__leaf_clk_i clknet_leaf_103_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_138_259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10610_ _05066_ memory\[50\]\[29\] _05203_ _05213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_25_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11590_ _05804_ _05805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__12693__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11496__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07311__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10541_ _05176_ _00311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_49_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_33_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13260_ _06831_ _02648_ _02650_ _02652_ _02653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_134_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10472_ _05064_ memory\[48\]\[28\] _05131_ _05140_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_118_clk_i clknet_5_23__leaf_clk_i clknet_leaf_118_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_40_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11768__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12211_ _06279_ _06416_ _06417_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_13191_ memory\[52\]\[24\] memory\[53\]\[24\] _06832_ _02585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_62_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_185_3929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12142_ memory\[60\]\[9\] memory\[61\]\[9\] _06273_ _06349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08142__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11567__I _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12073_ memory\[56\]\[8\] memory\[57\]\[8\] memory\[58\]\[8\] memory\[59\]\[8\] _06138_
+ _06280_ _06281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_60_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07981__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11024_ _05070_ memory\[56\]\[31\] _05398_ _05433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12599__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10923__I1 _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15832_ _00791_ clknet_leaf_134_clk_i memory\[9\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07780__I _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15763_ _00722_ clknet_leaf_133_clk_i memory\[62\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12825__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12975_ _05686_ _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11008__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10687__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14714_ _01753_ clknet_leaf_28_clk_i memory\[2\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11926_ memory\[62\]\[6\] memory\[63\]\[6\] _05868_ _06136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15694_ _00653_ clknet_leaf_255_clk_i memory\[60\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09701__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_169_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14645_ _01684_ clknet_leaf_80_clk_i memory\[27\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11857_ _06014_ _06036_ _06052_ _06068_ _06069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XTAP_TAPCELL_ROW_64_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13223__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_1066 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10439__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10808_ _05318_ _00436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14576_ _01615_ clknet_leaf_97_clk_i memory\[25\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13250__A1 _02167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_32_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11788_ memory\[62\]\[4\] memory\[63\]\[4\] _05868_ _06000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09500__I _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13527_ _05768_ _02911_ _02913_ _02915_ _02916_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_60_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_55_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10739_ _05058_ memory\[52\]\[25\] _05276_ _05282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13458_ memory\[12\]\[28\] memory\[13\]\[28\] _05769_ _02848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09057__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07020__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12409_ _06610_ _06612_ _06613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08804__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13389_ _02779_ _02780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_24_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09148__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15128_ _00087_ clknet_leaf_7_clk_i memory\[42\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08052__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_82_clk_i clknet_5_20__leaf_clk_i clknet_leaf_82_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11477__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07950_ _03206_ memory\[19\]\[26\] _03733_ _03740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15059_ _00018_ clknet_leaf_11_clk_i memory\[40\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_134_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08987__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06901_ net29 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_07881_ _03703_ _01204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_143_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09620_ _04672_ _01974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_97_clk_i clknet_5_20__leaf_clk_i clknet_leaf_97_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09780__I1 _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13069__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07791__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09551_ _04634_ _01943_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08502_ _04050_ _01478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09482_ _04587_ memory\[35\]\[6\] _04575_ _04588_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_188_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_176_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_20_clk_i clknet_5_5__leaf_clk_i clknet_leaf_20_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_148_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09611__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08433_ _03775_ memory\[20\]\[11\] _04012_ _04014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10757__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11940__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13241__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08364_ _03977_ _01413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09296__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08227__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07315_ memory\[11\]\[19\] _03348_ _03390_ _03400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_59_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_189_4007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_35_clk_i clknet_5_18__leaf_clk_i clknet_leaf_35_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_189_4018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08295_ _03772_ memory\[18\]\[10\] _03940_ _03941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10850__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08026__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_119_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07246_ _03358_ _00914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_6_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12771__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10492__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07177_ memory\[39\]\[1\] _03311_ _03309_ _03312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_446 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_41_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10602__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08897__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_855 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09220__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13308__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09818_ memory\[3\]\[24\] _03199_ _04773_ _04778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09749_ _04625_ memory\[38\]\[24\] _04736_ _04741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13155__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_336_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12760_ _02115_ _02130_ _02145_ _02160_ _02161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__13480__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11330__I1 _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11711_ _05914_ _05917_ _05920_ _05924_ _05925_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_68_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12946__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12691_ memory\[22\]\[16\] memory\[23\]\[16\] _06751_ _02093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10667__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_178_3799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11850__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_511 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14430_ _01469_ clknet_leaf_352_clk_i memory\[21\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11642_ _05856_ _05857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_154_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13232__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12167__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14361_ _01400_ clknet_leaf_106_clk_i memory\[18\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11573_ _05701_ _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_25_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput18 data_i[1] net18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13312_ memory\[62\]\[26\] memory\[63\]\[26\] _02448_ _02704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_64_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10524_ _05047_ memory\[4\]\[20\] _05167_ _05168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09039__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput29 data_i[2] net29 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10841__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14292_ _01331_ clknet_leaf_94_clk_i memory\[29\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13243_ _02358_ _02629_ _02636_ _02637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10455_ _05108_ _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_122_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13174_ _02568_ _02569_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_0_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10386_ _05094_ _00238_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12125_ memory\[30\]\[8\] memory\[31\]\[8\] _06193_ _06333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_176_Right_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_20_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08600__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12056_ _05788_ _06264_ _05792_ _06265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11007_ _05424_ _00529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15815_ _00774_ clknet_leaf_211_clk_i memory\[9\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_133_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15746_ _00705_ clknet_leaf_304_clk_i memory\[62\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12958_ _02209_ _02350_ _02353_ _02355_ _02356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07015__I net30 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13461__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11909_ _05918_ _06119_ _05775_ _06120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15677_ _00636_ clknet_leaf_336_clk_i memory\[60\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10577__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12889_ _06607_ _02287_ _02086_ _02288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_169_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_118_719 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14628_ _01667_ clknet_leaf_406_clk_i memory\[27\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_538 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_60_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14559_ _01598_ clknet_leaf_353_clk_i memory\[25\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_126_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07886__S _03697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07100_ _03267_ _03268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08080_ _03764_ memory\[15\]\[6\] _03819_ _03826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_3_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11880__S1 _06090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07031_ _03230_ _00827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_114_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_10_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_130_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_67_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11201__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_11_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_77_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_77_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08982_ _04319_ _01689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_285_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_143_Right_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_162_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07933_ _03181_ memory\[19\]\[18\] _03722_ _03731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13128__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12501__A3 _06702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07864_ _03694_ _01196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07764__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07126__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09603_ _04663_ _01966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07795_ _03178_ memory\[6\]\[17\] _03650_ _03658_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_27_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09534_ _03196_ _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_116_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09341__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09465_ _04576_ _01915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_4_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08416_ _03758_ memory\[20\]\[3\] _04001_ _04005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09269__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09396_ _04539_ _01883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_11_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11076__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08347_ _03968_ _01405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10286__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10823__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_116_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08278_ _03756_ memory\[18\]\[2\] _03929_ _03932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_34_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11871__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_134_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07229_ memory\[39\]\[18\] _03346_ _03330_ _03347_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10240_ _04637_ memory\[45\]\[30\] _04968_ _05002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09441__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11623__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10171_ _04965_ _00152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10950__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_110_Right_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09516__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08420__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13930_ _00969_ clknet_leaf_210_clk_i memory\[8\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_35_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06939__I _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07036__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_1225 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13861_ _00900_ clknet_leaf_404_clk_i memory\[39\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_83_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15600_ _00559_ clknet_leaf_176_clk_i memory\[57\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12812_ _02211_ _02212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_9_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13792_ _00831_ clknet_leaf_343_clk_i memory\[16\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12256__A2 _06460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09251__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11303__I1 _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15531_ _00490_ clknet_leaf_240_clk_i memory\[55\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12743_ _06318_ _02139_ _02141_ _02143_ _02144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__11580__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08180__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15462_ _00421_ clknet_leaf_299_clk_i memory\[53\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13205__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12674_ _06322_ _06873_ _06461_ _06874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_154_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14413_ _01452_ clknet_leaf_188_clk_i memory\[20\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11067__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11625_ _05732_ _05835_ _05837_ _05839_ _05840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_15393_ _00352_ clknet_leaf_327_clk_i memory\[51\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_13_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12803__I1 memory\[39\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11767__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13501__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14344_ _01383_ clknet_leaf_206_clk_i memory\[18\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11556_ _05681_ _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_25_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10507_ _05031_ memory\[4\]\[12\] _05156_ _05159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14275_ _01314_ clknet_leaf_355_clk_i memory\[29\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11487_ memory\[4\]\[0\] memory\[5\]\[0\] _05702_ _05703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13226_ _02216_ _02619_ _02620_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_0_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10438_ _05122_ _00262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_94_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09432__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12192__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11956__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10860__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13157_ _02337_ _02547_ _02549_ _02551_ _02552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_55_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10369_ _05029_ memory\[47\]\[11\] _05084_ _05086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_29_Left_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_55_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12108_ _05741_ _06315_ _06316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__09426__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08330__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13088_ _02337_ _02479_ _02481_ _02483_ _02484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_72_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_72_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12039_ _06247_ _06248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_40_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07746__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11691__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07580_ _03163_ memory\[0\]\[12\] _03541_ _03544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15729_ _00688_ clknet_leaf_162_clk_i memory\[61\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11490__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08171__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_38_Left_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_150_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09250_ _04461_ _01815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10100__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_138_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_141_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_150_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08201_ _03890_ _01337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_56_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09181_ _04241_ memory\[30\]\[28\] _04416_ _04425_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_84_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11758__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08132_ _03816_ memory\[15\]\[31\] _03818_ _03853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_79_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10805__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_55_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08505__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_79_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11853__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12535__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_151_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08063_ _03220_ _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XFILLER_0_183_1070 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13055__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07014_ _03216_ _00824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_105_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_47_Left_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_144_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11930__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_08965_ _04229_ memory\[27\]\[22\] _04308_ _04311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07916_ _03710_ _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08896_ _04274_ _01648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13683__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input24_I data_i[25] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07847_ _03685_ _01188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_07778_ _03153_ memory\[6\]\[9\] _03639_ _03649_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12089__I2 memory\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_56_Left_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_67_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09517_ _04611_ _01932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11614__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11997__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11106__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_175_3747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09448_ _04566_ _01908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11049__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_164_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09379_ _04235_ memory\[33\]\[25\] _04524_ _04530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11410_ _05615_ _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_10_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12390_ memory\[44\]\[12\] memory\[45\]\[12\] _06319_ _06594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_50_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09662__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_62_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_995 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11341_ _05601_ _00686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14060_ _01099_ clknet_leaf_214_clk_i memory\[10\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_1105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11272_ _05564_ _00654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_127_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13011_ memory\[14\]\[21\] memory\[15\]\[21\] _02193_ _02408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10223_ _04993_ _00176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08150__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10154_ _04619_ memory\[44\]\[21\] _04955_ _04957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11575__I _03113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14962_ _02001_ clknet_leaf_72_clk_i memory\[37\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_10__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10085_ _04920_ _00111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_50_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13913_ _00952_ clknet_leaf_134_clk_i memory\[11\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14893_ _01932_ clknet_leaf_51_clk_i memory\[35\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13844_ _00883_ clknet_leaf_114_clk_i memory\[13\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_18_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_175_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11524__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_18_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11288__I0 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13775_ _00814_ clknet_leaf_171_clk_i memory\[14\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_39 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10987_ _05033_ memory\[56\]\[13\] _05410_ _05414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_233_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11016__S _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11988__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12726_ memory\[8\]\[17\] memory\[9\]\[17\] memory\[10\]\[17\] memory\[11\]\[17\]
+ _06582_ _06721_ _02127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_15514_ _00473_ clknet_leaf_379_clk_i memory\[54\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07900__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15445_ _00404_ clknet_leaf_263_clk_i memory\[52\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12657_ memory\[14\]\[16\] memory\[15\]\[16\] _06302_ _06857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13231__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_5_19__f_clk_i clknet_2_2_0_clk_i clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_25_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11608_ memory\[0\]\[1\] memory\[1\]\[1\] memory\[2\]\[1\] memory\[3\]\[1\] _05711_
+ _03748_ _05823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_155_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_96_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15376_ _00335_ clknet_leaf_157_clk_i memory\[50\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12588_ _06713_ _06784_ _06786_ _06788_ _06789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_68_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_96_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12355__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14327_ _01366_ clknet_leaf_115_clk_i memory\[17\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10412__A1 _03227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11539_ memory\[46\]\[0\] memory\[47\]\[0\] _05754_ _05755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_399 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_57_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14258_ _01297_ clknet_leaf_114_clk_i memory\[15\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09405__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13588__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11686__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13209_ _05772_ _02602_ _02195_ _02603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11212__I0 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14189_ _01228_ clknet_leaf_194_clk_i memory\[19\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11912__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07963__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09156__S _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11485__I _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08750_ net74 _03855_ _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_174_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08995__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07719__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12012__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13665__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07701_ _03608_ _01119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08681_ net73 _03855_ _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_75_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08392__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07195__I1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_139_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07632_ _03138_ memory\[10\]\[4\] _03567_ _03572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_109_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12310__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13417__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08794__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07404__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07563_ _03138_ memory\[0\]\[4\] _03530_ _03535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08144__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11979__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_441_clk_i clknet_5_1__leaf_clk_i clknet_leaf_441_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09302_ _04489_ _01839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_192_4058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_192_4069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07494_ memory\[59\]\[4\] _03317_ _03493_ _03498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07203__I _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09892__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_61_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_63_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_153_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09233_ _04224_ memory\[31\]\[20\] _04452_ _04453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10765__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_748 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_111_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09164_ _04393_ _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_90_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08235__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12265__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08115_ _03844_ _01297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_47_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09095_ _04379_ _01742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_131_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_435_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13028__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_131_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08046_ _03804_ memory\[12\]\[25\] _03794_ _03805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_47_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11596__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12156__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11203__I0 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11903__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07958__I0 _03218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13096__B _02489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09997_ _04598_ memory\[42\]\[11\] _04872_ _04874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_182_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08948_ _04212_ memory\[27\]\[14\] _04297_ _04302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10005__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_129_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08879_ _04265_ _01640_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_4_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_70 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07186__I1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10910_ memory\[55\]\[9\] _03152_ _05363_ _05373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10190__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11890_ _05699_ _06093_ _06100_ _06101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_98_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_19_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_98_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10841_ _05024_ memory\[54\]\[9\] _05326_ _05336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13503__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11809__I2 memory\[2\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_409_clk_i clknet_5_2__leaf_clk_i clknet_leaf_409_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_15_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13560_ _02948_ net61 _02382_ _02949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10772_ _05299_ _00419_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12511_ _05675_ _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
X_13491_ _02371_ _02880_ _02373_ _02881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12954__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10675__S _05240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15230_ _00189_ clknet_leaf_416_clk_i memory\[46\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_136_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12442_ _06162_ _06644_ _06645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_81_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09635__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_151_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12175__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15161_ _00120_ clknet_leaf_3_clk_i memory\[43\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12373_ _06155_ _06572_ _06574_ _06576_ _06577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12490__S1 _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07984__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14112_ _01151_ clknet_leaf_308_clk_i memory\[6\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11324_ memory\[61\]\[11\] _03159_ _05591_ _05593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15092_ _00051_ clknet_leaf_11_clk_i memory\[41\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12147__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14043_ _01082_ clknet_leaf_395_clk_i memory\[0\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11255_ _03332_ memory\[60\]\[11\] _05554_ _05556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_52_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10206_ _04984_ _00168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11186_ _05519_ _00613_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10137_ _04602_ memory\[44\]\[13\] _04944_ _04948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_13_Right_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14945_ _01984_ clknet_leaf_437_clk_i memory\[37\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10068_ _04911_ _00103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07177__I1 _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12130__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14876_ _01915_ clknet_leaf_425_clk_i memory\[35\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09503__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13827_ _00866_ clknet_leaf_284_clk_i memory\[13\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08126__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_384_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13758_ _00797_ clknet_leaf_280_clk_i memory\[14\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_85_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08677__I1 _03371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07023__I net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12709_ memory\[54\]\[17\] memory\[55\]\[17\] _06421_ _02110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10484__I1 memory\[4\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10585__S _05192_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13689_ _03074_ _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13258__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15428_ _00387_ clknet_leaf_316_clk_i memory\[52\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08055__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Right_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_14_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12386__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11433__I0 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15359_ _00318_ clknet_leaf_348_clk_i memory\[50\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_13_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12138__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09920_ _04589_ memory\[41\]\[7\] _04825_ _04833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12305__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09851_ _04796_ _00001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08802_ _04217_ _01611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09782_ memory\[3\]\[7\] _03146_ _04751_ _04759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06994_ _03201_ _00819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_31_Right_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13638__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_146_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08733_ _03802_ memory\[24\]\[24\] _04168_ _04173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08365__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13136__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08664_ _04136_ _01554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12040__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_1_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10172__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07134__S _03279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07615_ _03215_ memory\[0\]\[29\] _03552_ _03562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_380_clk_i clknet_5_12__leaf_clk_i clknet_leaf_380_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_117_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08595_ _04099_ _01522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08029__I _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07546_ memory\[59\]\[29\] _03369_ _03515_ _03525_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_129_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07477_ _03487_ _01016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_40_Right_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_147_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07340__I1 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09216_ _04208_ memory\[31\]\[12\] _04441_ _04444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_395_clk_i clknet_5_6__leaf_clk_i clknet_leaf_395_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_106_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09617__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12377__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09147_ _04407_ _01766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_32_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_20_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09078_ _04206_ memory\[2\]\[11\] _04369_ _04371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12129__A1 _05914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08029_ _03186_ _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_187_3971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07309__S _03390_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11040_ _05018_ memory\[57\]\[6\] _05435_ _05442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_333_clk_i clknet_5_8__leaf_clk_i clknet_leaf_333_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_output55_I net55 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13554__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12991_ memory\[56\]\[21\] memory\[57\]\[21\] memory\[58\]\[21\] memory\[59\]\[21\]
+ _06827_ _02171_ _02388_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08356__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12301__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1030 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14730_ _01769_ clknet_leaf_131_clk_i memory\[30\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11942_ _06149_ _06151_ _06152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06947__I _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07044__S _03229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_348_clk_i clknet_5_8__leaf_clk_i clknet_leaf_348_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_87_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_1059 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14661_ _01700_ clknet_leaf_360_clk_i memory\[28\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11873_ _05676_ _06079_ _06081_ _06083_ _06084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_129_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13612_ _02501_ _02999_ _03000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_131_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10824_ _05327_ _00443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14592_ _01631_ clknet_leaf_415_clk_i memory\[26\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08659__I1 _03353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09856__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12684__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13543_ _02336_ _02924_ _02931_ _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_94_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10755_ _05004_ memory\[53\]\[0\] _05290_ _05291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_45_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13474_ _02863_ _02864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_192_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10686_ _05253_ _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_62_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15213_ _00172_ clknet_leaf_386_clk_i memory\[45\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11415__I0 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12425_ _06276_ _06627_ _06001_ _06628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_23_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12463__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15144_ _00103_ clknet_leaf_29_clk_i memory\[43\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12356_ memory\[56\]\[12\] memory\[57\]\[12\] memory\[58\]\[12\] memory\[59\]\[12\]
+ _06138_ _06280_ _06560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_105_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_306 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11307_ memory\[61\]\[3\] _03134_ _05580_ _05584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_10_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15075_ _00034_ clknet_leaf_433_clk_i memory\[41\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12125__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12287_ _06492_ _00741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14026_ _01065_ clknet_leaf_218_clk_i memory\[0\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11238_ _03315_ memory\[60\]\[3\] _05543_ _05547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11964__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11169_ _05510_ _00605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09434__S _04549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10154__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14928_ _01967_ clknet_leaf_67_clk_i memory\[36\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_141_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14859_ _01898_ clknet_leaf_53_clk_i memory\[34\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07400_ _03209_ memory\[8\]\[27\] _03437_ _03445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_102_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08380_ _03985_ _01421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_102_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_130_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07331_ _03408_ _00949_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_441 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__I1 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07262_ _03214_ _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_171_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_182_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09001_ _04197_ memory\[28\]\[7\] _04322_ _04330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11406__I0 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_472 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07193_ _03322_ _00897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13651__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07086__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09609__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08513__S _04048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12543__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_148_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09903_ _04823_ _00026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_165_3554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09834_ _03113_ _03304_ _04786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__06968__S _03157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_55_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_126_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09765_ _03376_ _03528_ _04749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_06977_ _03187_ memory\[14\]\[20\] _03188_ _03189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08338__I0 _03816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08716_ _03785_ memory\[24\]\[16\] _04157_ _04164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09696_ _04712_ _02010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10145__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09143__I _04393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08647_ _04127_ _01546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10289__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07799__S _03650_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08578_ _04090_ _01514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09838__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12718__B _06707_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07529_ _03516_ _01039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11622__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12693__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07313__I1 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11114__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_783 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_106_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10540_ _05064_ memory\[4\]\[28\] _05167_ _05176_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_729 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10471_ _05139_ _00278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_157_Right_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_40_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12210_ memory\[56\]\[10\] memory\[57\]\[10\] memory\[58\]\[10\] memory\[59\]\[10\]
+ _06138_ _06280_ _06416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09519__S _04596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13190_ _02163_ _02579_ _02581_ _02583_ _02584_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_60_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_680 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_332_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12141_ _06348_ _00739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_341 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1090 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_12072_ _03116_ _06280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xclkbuf_leaf_272_clk_i clknet_5_13__leaf_clk_i clknet_leaf_272_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_102_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08577__I0 _03783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12522__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11784__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11023_ _05432_ _00537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15831_ _00790_ clknet_leaf_129_clk_i memory\[9\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_287_clk_i clknet_5_15__leaf_clk_i clknet_leaf_287_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_86_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12974_ memory\[22\]\[20\] memory\[23\]\[20\] _06751_ _02372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15762_ _00721_ clknet_leaf_178_clk_i memory\[62\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07001__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14713_ _01752_ clknet_leaf_59_clk_i memory\[2\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11925_ _06134_ _06135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_169_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_47_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_1_clk_i clknet_5_4__leaf_clk_i clknet_leaf_1_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15693_ _00652_ clknet_leaf_236_clk_i memory\[60\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_840 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_210_clk_i clknet_5_30__leaf_clk_i clknet_leaf_210_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14644_ _01683_ clknet_leaf_95_clk_i memory\[27\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08892__I _04249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11856_ _05767_ _06059_ _06067_ _06068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_64_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_158 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12589__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07502__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10807_ _05058_ memory\[53\]\[25\] _05312_ _05318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14575_ _01614_ clknet_leaf_125_clk_i memory\[25\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11787_ _05998_ _05999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_32_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08501__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11024__S _05398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13526_ _05777_ _02914_ _02915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_TAPCELL_ROW_60_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10738_ _05281_ _00403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_125_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_770 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_225_clk_i clknet_5_27__leaf_clk_i clknet_leaf_225_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13457_ _05747_ _02842_ _02844_ _02846_ _02847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_82_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10669_ memory\[51\]\[24\] _03199_ _05240_ _05245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_124_Right_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_153_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12408_ memory\[24\]\[12\] memory\[25\]\[12\] memory\[26\]\[12\] memory\[27\]\[12\]
+ _06472_ _06611_ _06612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_88_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_639 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13388_ memory\[4\]\[27\] memory\[5\]\[27\] _05789_ _02779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12339_ _05914_ _06539_ _06541_ _06543_ _06544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_15127_ _00086_ clknet_leaf_10_clk_i memory\[42\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_10_Left_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_121_683 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15058_ _00017_ clknet_leaf_13_clk_i memory\[40\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_120_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11694__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06900_ _03130_ _00796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14009_ _01048_ clknet_leaf_268_clk_i memory\[59\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07880_ _03203_ memory\[7\]\[25\] _03697_ _03703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10375__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07971__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13194__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13069__A2 _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09550_ _04633_ memory\[35\]\[28\] _04617_ _04634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_160_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08501_ _03775_ memory\[21\]\[11\] _04048_ _04050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09481_ _03143_ _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__11875__I0 memory\[4\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_144_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08432_ _04013_ _01445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_281_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08363_ _03772_ memory\[1\]\[10\] _03976_ _03977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07314_ _03399_ _00941_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_22_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_189_4008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08294_ _03928_ _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_34_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11869__S _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07245_ memory\[39\]\[23\] _03357_ _03351_ _03358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10773__S _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07059__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09339__S _04502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__08243__S _03904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07176_ _03128_ _03311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_15_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08042__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_180_3838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09817_ _04777_ _02066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10013__S _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10118__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09748_ _04740_ _02034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12363__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10669__I1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10948__S _05385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09679_ _04623_ memory\[37\]\[23\] _04700_ _04704_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08731__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07534__I1 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11710_ _05921_ _05923_ _05924_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_166_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12690_ _02091_ _02092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08418__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07322__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11641_ memory\[20\]\[1\] memory\[21\]\[1\] _05785_ _05856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14360_ _01399_ clknet_leaf_106_clk_i memory\[18\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_64_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11572_ _05752_ _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_0_65_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07121__I _03267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13311_ _02702_ _02703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10523_ _05144_ _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
Xinput19 data_i[20] net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_14291_ _01330_ clknet_leaf_83_clk_i memory\[29\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10683__S _05217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13242_ _02367_ _02631_ _02633_ _02635_ _02636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__09249__S _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10454_ _05130_ _00270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08798__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11578__I _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12743__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13173_ memory\[20\]\[23\] memory\[21\]\[23\] _02368_ _02568_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10385_ _05045_ memory\[47\]\[19\] _05084_ _05094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12124_ _06331_ _06332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_27_1299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11929__S0 _06138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12055_ memory\[22\]\[7\] memory\[23\]\[7\] _06062_ _06264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11006_ _05052_ memory\[56\]\[22\] _05421_ _05424_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_189_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15814_ _00773_ clknet_leaf_216_clk_i memory\[9\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_29_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15745_ _00704_ clknet_leaf_305_clk_i memory\[62\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_133_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12957_ _02216_ _02354_ _02355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10858__S _05337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_59_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08722__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07525__I1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11482__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11908_ memory\[30\]\[5\] memory\[31\]\[5\] _05773_ _06119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08328__S _03951_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15676_ _00635_ clknet_leaf_335_clk_i memory\[60\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12888_ memory\[30\]\[19\] memory\[31\]\[19\] _02084_ _02287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14627_ _01666_ clknet_leaf_413_clk_i memory\[27\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11839_ _05748_ _06046_ _06048_ _06050_ _06051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_28_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_164_clk_i clknet_5_25__leaf_clk_i clknet_leaf_164_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_126_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14558_ _01597_ clknet_leaf_415_clk_i memory\[25\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_3_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12982__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13509_ _05719_ _02897_ _05739_ _02898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14489_ _01528_ clknet_leaf_106_clk_i memory\[22\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_148_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07030_ _03111_ memory\[16\]\[0\] _03229_ _03230_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08789__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_179_clk_i clknet_5_28__leaf_clk_i clknet_leaf_179_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_23_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10596__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_2_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_77_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_114_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_228_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08981_ _04245_ memory\[27\]\[30\] _04285_ _04319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_139_64 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07932_ _03730_ _01228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_102_clk_i clknet_5_21__leaf_clk_i clknet_leaf_102_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_162_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08797__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10348__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07863_ _03178_ memory\[7\]\[17\] _03686_ _03694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08961__I0 _04224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09602_ _04614_ memory\[36\]\[19\] _04653_ _04663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_155_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07794_ _03657_ _01163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_117_clk_i clknet_5_23__leaf_clk_i clknet_leaf_117_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09533_ _04622_ _01937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09464_ _04573_ memory\[35\]\[0\] _04575_ _04576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwire76 _03266_ net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_93_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08415_ _04004_ _01437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_8_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09395_ _04181_ memory\[34\]\[0\] _04538_ _04539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08346_ _03756_ memory\[1\]\[2\] _03965_ _03968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_184_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__06981__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_7_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_173_3697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_11_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08277_ _03931_ _01372_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_190_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_172_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_751 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__S _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07228_ _03180_ _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_104_425 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_134_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_134_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12725__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07159_ _03212_ memory\[13\]\[28\] _03290_ _03299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10587__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10170_ _04635_ memory\[44\]\[29\] _04955_ _04965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08701__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13319__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10339__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12223__S _06156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13150__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13860_ _00899_ clknet_leaf_396_clk_i memory\[39\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_83_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09532__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12811_ memory\[44\]\[18\] memory\[45\]\[18\] _02210_ _02211_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13791_ _00830_ clknet_leaf_365_clk_i memory\[16\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08704__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07507__I1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15530_ _00489_ clknet_leaf_242_clk_i memory\[55\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06955__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12742_ _06325_ _02142_ _02143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__08148__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10511__I0 _05035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_81_clk_i clknet_5_20__leaf_clk_i clknet_leaf_81_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_69_Right_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12893__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15461_ _00420_ clknet_leaf_317_clk_i memory\[53\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12673_ memory\[46\]\[16\] memory\[47\]\[16\] _06596_ _06873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_388 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07987__S _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14412_ _01451_ clknet_leaf_192_clk_i memory\[20\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11624_ _05741_ _05838_ _05839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_155_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_177_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15392_ _00351_ clknet_leaf_334_clk_i memory\[51\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_182_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_526 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_13_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_53_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12964__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14343_ _01382_ clknet_leaf_205_clk_i memory\[18\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_53_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11555_ _05770_ _05771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_96_clk_i clknet_5_20__leaf_clk_i clknet_leaf_96_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_163_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10506_ _05158_ _00294_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14274_ _01313_ clknet_leaf_408_clk_i memory\[29\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11486_ _05701_ _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_123_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13225_ memory\[40\]\[24\] memory\[41\]\[24\] memory\[42\]\[24\] memory\[43\]\[24\]
+ _06875_ _02217_ _02619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_111_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10437_ _05029_ memory\[48\]\[11\] _05120_ _05122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_94_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09707__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_78_Right_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_110_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13156_ _02344_ _02550_ _02551_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10368_ _05085_ _00229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_55_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13229__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12107_ memory\[32\]\[8\] memory\[33\]\[8\] memory\[34\]\[8\] memory\[35\]\[8\] _06314_
+ _05743_ _06315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_97_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13087_ _02344_ _02482_ _02483_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10299_ _05041_ memory\[46\]\[17\] _05027_ _05042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13141__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09506__I _03168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12038_ memory\[44\]\[7\] memory\[45\]\[7\] _05749_ _06247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_72_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_34_clk_i clknet_5_7__leaf_clk_i clknet_leaf_34_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11972__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07026__I _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_178_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13989_ _01028_ clknet_leaf_318_clk_i memory\[59\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_177_428 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_87_Right_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15728_ _00687_ clknet_leaf_147_clk_i memory\[61\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08058__S _03794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_49_clk_i clknet_5_18__leaf_clk_i clknet_leaf_49_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12088__B _06018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10387__I _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_138_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15659_ _00618_ clknet_leaf_244_clk_i memory\[5\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_138_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_118_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08200_ _03814_ memory\[29\]\[30\] _03856_ _03890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09180_ _04424_ _01782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06882__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_69_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08131_ _03852_ _01305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_173_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_79_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_172_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11212__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07682__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08062_ _03815_ _01273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_183_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13055__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_71_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07013_ _03215_ memory\[14\]\[29\] _03188_ _03216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_96_Right_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_102_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09617__S _04664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_379_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12551__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11946__I _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08964_ _04310_ _01680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_45_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09187__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07915_ _03721_ _01220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08895_ _04227_ memory\[26\]\[21\] _04272_ _04274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07846_ _03153_ memory\[7\]\[9\] _03675_ _03685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10741__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09352__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input17_I data_i[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_431_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_116_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10498__S _05145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07777_ _03648_ _01155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12238__A3 _06443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_3_Left_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_155_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09516_ _04610_ memory\[35\]\[17\] _04596_ _04611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09447_ _04235_ memory\[34\]\[25\] _04560_ _04566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_176_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_175_3748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_137_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_137_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09378_ _04529_ _01875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09111__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08329_ _03958_ _01397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_10_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_380 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11340_ memory\[61\]\[19\] _03183_ _05591_ _05601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13746__I0 _03365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11271_ _03348_ memory\[60\]\[19\] _05554_ _05564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13010_ _02406_ _02407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_132_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10222_ _04619_ memory\[45\]\[21\] _04991_ _04993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11921__A2 _06101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10153_ _04956_ _00143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09326__I _04501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10084_ _04616_ memory\[43\]\[20\] _04919_ _04920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14961_ _02000_ clknet_leaf_18_clk_i memory\[37\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12888__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08925__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13912_ _00951_ clknet_leaf_134_clk_i memory\[11\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14892_ _01931_ clknet_leaf_52_clk_i memory\[35\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_57_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13843_ _00882_ clknet_leaf_117_clk_i memory\[13\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_97_551 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10201__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13774_ _00813_ clknet_leaf_173_clk_i memory\[14\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10986_ _05413_ _00519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_168_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09350__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15513_ _00472_ clknet_leaf_385_clk_i memory\[54\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12725_ _06717_ _02125_ _06304_ _02126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_15444_ _00403_ clknet_leaf_262_clk_i memory\[52\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08606__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12656_ _06855_ _06856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_127_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_824 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12937__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1044 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11607_ _05705_ _05821_ _05708_ _05822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12587_ _06720_ _06787_ _06788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_25_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15375_ _00334_ clknet_leaf_256_clk_i memory\[50\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_96_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10799__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11032__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_170_648 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14326_ _01365_ clknet_leaf_111_clk_i memory\[17\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10412__A2 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11538_ _05701_ _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_41_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14257_ _01296_ clknet_leaf_114_clk_i memory\[15\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11469_ memory\[54\]\[0\] memory\[55\]\[0\] _05684_ _05685_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10871__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09437__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13208_ memory\[14\]\[24\] memory\[15\]\[24\] _02193_ _02602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_380_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14188_ _01227_ clknet_leaf_192_clk_i memory\[19\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10176__A1 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13139_ _06848_ _02533_ _06707_ _02534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09169__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input9_I data_i[11] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07700_ _03138_ memory\[63\]\[4\] _03603_ _03608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08680_ _04144_ _01562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_139_1168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07631_ _03571_ _01086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_109_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11715__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07562_ _03534_ _01054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_49_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09341__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09301_ _04224_ memory\[32\]\[20\] _04488_ _04489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09900__S _04788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_192_4059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07493_ _03497_ _01022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_76_757 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_174_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09232_ _04429_ _04452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_57_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07420__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12928__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09163_ _04415_ _01774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11450__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12038__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_1098 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_170_3656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08114_ _03798_ memory\[15\]\[22\] _03841_ _03844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07655__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_659 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08315__I _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09094_ _04222_ memory\[2\]\[19\] _04369_ _04379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_473 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_131_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_1236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13028__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11877__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08045_ _03202_ _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_114_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12156__A2 _06355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13353__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08080__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_125_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10962__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09996_ _04873_ _00069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_792 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08947_ _04301_ _01672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_129_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08907__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11667__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08878_ _04210_ memory\[26\]\[13\] _04261_ _04265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10714__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09082__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_4_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_19_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_4_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07829_ _03676_ _01179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11117__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10840_ _05335_ _00451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09810__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_15_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12711__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10771_ _05022_ memory\[53\]\[8\] _05290_ _05299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10956__S _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13332__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12510_ _06155_ _06705_ _06708_ _06711_ _06712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_137_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13490_ memory\[22\]\[28\] memory\[23\]\[28\] _05754_ _02880_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08426__S _04001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07330__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12919__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12441_ memory\[0\]\[13\] memory\[1\]\[13\] memory\[2\]\[13\] memory\[3\]\[13\] _06020_
+ _06090_ _06644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_47_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12372_ _06162_ _06575_ _06576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_129_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15160_ _00119_ clknet_leaf_7_clk_i memory\[43\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_65_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13719__I0 _03338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14111_ _01150_ clknet_leaf_285_clk_i memory\[6\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_105_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11323_ _05592_ _00677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12970__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10691__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07271__A1 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15091_ _00050_ clknet_leaf_11_clk_i memory\[41\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09399__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14042_ _01081_ clknet_leaf_395_clk_i memory\[0\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11254_ _05555_ _00645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08161__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13287__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11586__I _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10205_ _04602_ memory\[45\]\[13\] _04980_ _04984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_52_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11185_ _03329_ memory\[5\]\[10\] _05518_ _05519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10136_ _04947_ _00135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_140_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12411__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11658__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14944_ _01983_ clknet_leaf_437_clk_i memory\[37\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10067_ _04600_ memory\[43\]\[12\] _04908_ _04911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10705__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09571__I0 _04583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14875_ _01914_ clknet_leaf_1_clk_i memory\[34\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12870__A3 _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13826_ _00865_ clknet_leaf_283_clk_i memory\[13\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_327_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09323__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09720__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12083__A1 _06142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_134_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13757_ _00796_ clknet_leaf_276_clk_i memory\[14\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10969_ _05404_ _00511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12708_ _02108_ _02109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_39_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08336__S _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13688_ _03115_ net75 _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_171_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13258__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_75_Left_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_183_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15427_ _00386_ clknet_leaf_315_clk_i memory\[52\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_54_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12639_ _05693_ _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_109_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13583__A1 _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15358_ _00317_ clknet_leaf_348_clk_i memory\[50\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_40_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_103_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14309_ _01348_ clknet_leaf_368_clk_i memory\[17\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_79_8 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15289_ _00248_ clknet_leaf_385_clk_i memory\[47\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07974__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13335__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09167__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1280 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11197__I0 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11897__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09850_ _04587_ memory\[40\]\[6\] _04789_ _04796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10106__S _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08801_ _04216_ memory\[25\]\[16\] _04204_ _04217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_84_Left_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_06993_ _03200_ memory\[14\]\[24\] _03188_ _03201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09781_ _04758_ _02049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08732_ _04172_ _01586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08663_ memory\[23\]\[23\] _03357_ _04132_ _04136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12161__I2 memory\[2\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_124_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07614_ _03561_ _01079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08594_ _03800_ memory\[22\]\[23\] _04095_ _04099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_191_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12074__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07545_ _03524_ _01047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_138_Right_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10776__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11121__I0 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_14_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_93_Left_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_118_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07876__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_431 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07476_ memory\[49\]\[29\] _03369_ _03477_ _03487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09215_ _04443_ _01798_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_51_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_401 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09146_ _04206_ memory\[30\]\[11\] _04405_ _04407_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13574__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07628__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08045__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09077_ _04370_ _01733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_20_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11680__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11400__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_4_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08028_ _03792_ _01262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_187_3972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11888__A1 _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10016__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_276_clk_i_I clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09805__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09979_ _04864_ _00061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13327__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12231__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12990_ _02167_ _02386_ _06690_ _02387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_98_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output48_I net48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09604__I _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09553__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_157_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11941_ memory\[48\]\[6\] memory\[49\]\[6\] memory\[50\]\[6\] memory\[51\]\[6\] _06010_
+ _06150_ _06151_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_170_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_98_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14660_ _01699_ clknet_leaf_361_clk_i memory\[28\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_169_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11872_ _05690_ _06082_ _06083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_169_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09305__I0 _04229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13611_ memory\[24\]\[30\] memory\[25\]\[30\] memory\[26\]\[30\] memory\[27\]\[30\]
+ _05742_ _02502_ _02999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12965__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10823_ _05004_ memory\[54\]\[0\] _05326_ _05327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14591_ _01630_ clknet_leaf_415_clk_i memory\[26\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11112__I0 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_105_Right_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_184_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06963__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07867__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13542_ _05676_ _02926_ _02928_ _02930_ _02931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__08156__S _03857_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10754_ _05289_ _05290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_153_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10685_ _03451_ _03750_ _05253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_13473_ memory\[44\]\[28\] memory\[45\]\[28\] _05678_ _02863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_35_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_63_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13565__A1 _05705_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15212_ _00171_ clknet_leaf_37_clk_i memory\[45\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_164_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12424_ memory\[62\]\[13\] memory\[63\]\[13\] _06557_ _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07619__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15143_ _00102_ clknet_leaf_22_clk_i memory\[43\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_129_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08292__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12355_ _06276_ _06558_ _06001_ _06559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_51_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11306_ _05583_ _00669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15074_ _00033_ clknet_leaf_442_clk_i memory\[41\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12286_ _06490_ net41 _06491_ _06492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14025_ _01064_ clknet_leaf_248_clk_i memory\[0\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11237_ _05546_ _00637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12205__I _03450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_440_clk_i clknet_5_0__leaf_clk_i clknet_leaf_440_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09715__S _04714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11168_ _03313_ memory\[5\]\[2\] _05507_ _05510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10119_ _04938_ _00127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11099_ _05473_ _00572_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_1086 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09544__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14927_ _01966_ clknet_leaf_65_clk_i memory\[36\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_320 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14858_ _01897_ clknet_leaf_45_clk_i memory\[34\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13809_ _00848_ clknet_leaf_117_clk_i memory\[16\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12056__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_102_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10596__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14789_ _01828_ clknet_leaf_401_clk_i memory\[32\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_86_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07330_ memory\[11\]\[26\] _03363_ _03401_ _03408_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_420 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_82_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_133_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_2_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07483__A1 _03376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07261_ _03368_ _00919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_412 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09000_ _04329_ _01697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13556__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13700__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07192_ memory\[39\]\[6\] _03321_ _03309_ _03322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_5_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13651__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11220__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10090__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_408_clk_i clknet_5_3__leaf_clk_i clknet_leaf_408_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09902_ _04639_ memory\[40\]\[31\] _04788_ _04823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_165_3544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_6_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09625__S _04641_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_09833_ _04785_ _02074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_126_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09764_ _04748_ _02042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06976_ _03125_ _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07145__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09535__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08715_ _04163_ _01578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_154_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09695_ _04639_ memory\[37\]\[31\] _04677_ _04712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08646_ memory\[23\]\[15\] _03340_ _04121_ _04127_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09360__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08577_ _03783_ memory\[22\]\[15\] _04084_ _04090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_138_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07528_ memory\[59\]\[20\] _03350_ _03515_ _03516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07849__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_0__f_clk_i clknet_2_0_0_clk_i clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_77_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07459_ _03478_ _01007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13547__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_49_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10470_ _05062_ memory\[48\]\[27\] _05131_ _05139_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08704__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_40_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09129_ _04189_ memory\[30\]\[3\] _04394_ _04398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_40_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08274__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12226__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_890 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12140_ _06347_ net70 _05802_ _06348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10081__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12071_ _05667_ _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_11022_ _05068_ memory\[56\]\[30\] _05398_ _05432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09535__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13565__B _05756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15830_ _00789_ clknet_leaf_134_clk_i memory\[9\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06958__I net14 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07055__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09526__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15761_ _00720_ clknet_leaf_178_clk_i memory\[62\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12973_ _05752_ _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_86_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14712_ _01751_ clknet_leaf_59_clk_i memory\[2\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11924_ memory\[60\]\[6\] memory\[61\]\[6\] _05656_ _06134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15692_ _00651_ clknet_leaf_222_clk_i memory\[60\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_47_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14643_ _01682_ clknet_leaf_96_clk_i memory\[27\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_386 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11855_ _05783_ _06061_ _06064_ _06066_ _06067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_184_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11305__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10806_ _05317_ _00435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14574_ _01613_ clknet_leaf_126_clk_i memory\[25\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_71_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11786_ memory\[60\]\[4\] memory\[61\]\[4\] _05656_ _05998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_172_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13525_ memory\[8\]\[29\] memory\[9\]\[29\] memory\[10\]\[29\] memory\[11\]\[29\]
+ _02473_ _05779_ _02914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_153_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_32_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10737_ _05056_ memory\[52\]\[24\] _05276_ _05281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_67_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13456_ _05759_ _02845_ _02846_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10668_ _05244_ _00370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_149_Left_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12407_ _03747_ _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_125_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10599_ _05207_ _00338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13387_ _02302_ _02770_ _02777_ _02778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__11040__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09509__I _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15126_ _00085_ clknet_leaf_6_clk_i memory\[42\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12338_ _05921_ _06542_ _06543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_2_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_1251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15057_ _00016_ clknet_leaf_16_clk_i memory\[40\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12269_ _05914_ _06469_ _06471_ _06474_ _06475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_121_695 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07029__I _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14008_ _01047_ clknet_leaf_266_clk_i memory\[59\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09445__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_143_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_394_clk_i clknet_5_6__leaf_clk_i clknet_leaf_394_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_170_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_158_Left_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12277__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_160_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_179_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08500_ _04049_ _01477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09480_ _04586_ _01920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_121_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_176_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_504 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08431_ _03772_ memory\[20\]\[10\] _04012_ _04013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12029__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_224_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08362_ _03964_ _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_86_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13321__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07313_ memory\[11\]\[18\] _03346_ _03390_ _03399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_22_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_22_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08293_ _03939_ _01380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_50_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_332_clk_i clknet_5_8__leaf_clk_i clknet_leaf_332_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_189_4009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_167_Left_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_61_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07244_ _03196_ _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_160_97 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_1020 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08524__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_119_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_5_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_119_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11949__I _05659_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08256__I0 _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07175_ _03310_ _00891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12201__A1 _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12046__S _05915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10063__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_347_clk_i clknet_5_8__leaf_clk_i clknet_leaf_347_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_112_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11885__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_100_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_EDGE_ROW_176_Left_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_180_3839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09816_ memory\[3\]\[23\] _03196_ _04773_ _04777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_185_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_154_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12268__A1 _05921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09747_ _04623_ memory\[38\]\[23\] _04736_ _04740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06959_ _03174_ _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_69_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12363__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_190_Right_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_90_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09678_ _04703_ _02001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_958 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09090__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07603__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08629_ memory\[23\]\[7\] _03323_ _04110_ _04118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_90_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11125__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11640_ _05768_ _05850_ _05852_ _05854_ _05855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_37_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12440__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10964__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11571_ _05786_ _05787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_135_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_505 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13340__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13310_ memory\[60\]\[26\] memory\[61\]\[26\] _02164_ _02702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10522_ _05166_ _00302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14290_ _01329_ clknet_leaf_82_clk_i memory\[29\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13241_ _02375_ _02634_ _02635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_126_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10453_ _05045_ memory\[48\]\[19\] _05120_ _05130_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_426_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10054__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09995__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13172_ _02494_ _02562_ _02564_ _02566_ _02567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_10384_ _05093_ _00237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12123_ memory\[28\]\[8\] memory\[29\]\[8\] _05915_ _06331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07470__I1 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09747__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12054_ _06262_ _06263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__11929__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13295__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_173_clk_i_I clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11005_ _05423_ _00528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15813_ _00772_ clknet_leaf_298_clk_i memory\[9\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12259__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06981__I0 _03191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15744_ _00703_ clknet_leaf_306_clk_i memory\[62\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_172_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12956_ memory\[40\]\[20\] memory\[41\]\[20\] memory\[42\]\[20\] memory\[43\]\[20\]
+ _06875_ _02217_ _02354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_88_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07513__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11907_ _06117_ _06118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_15675_ _00634_ clknet_leaf_396_clk_i memory\[5\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12887_ _02285_ _02286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_74_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13303__S0 _02233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14626_ _01665_ clknet_leaf_409_clk_i memory\[27\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11838_ _05760_ _06049_ _06050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_23_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08486__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14557_ _01596_ clknet_leaf_407_clk_i memory\[25\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11769_ _05981_ _05982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10293__I0 _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13508_ memory\[54\]\[29\] memory\[55\]\[29\] _02312_ _02897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08344__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_98_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14488_ _01527_ clknet_leaf_109_clk_i memory\[22\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13439_ _05705_ _02828_ _05756_ _02829_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_144_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_84_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09986__I0 _04587_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_77_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15109_ _00068_ clknet_leaf_445_clk_i memory\[42\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_41_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08980_ _04318_ _01688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_121_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09175__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09738__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07931_ _03178_ memory\[19\]\[17\] _03722_ _03730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_162_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12042__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08410__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07862_ _03693_ _01195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10114__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09601_ _04662_ _01965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07793_ _03175_ memory\[6\]\[16\] _03650_ _03657_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06972__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13425__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09532_ _04621_ memory\[35\]\[22\] _04617_ _04622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_91_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_189_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09910__I0 _04579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09463_ _04574_ _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_148_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_375_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08414_ _03756_ memory\[20\]\[2\] _04001_ _04004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09394_ _04537_ _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_65_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_191_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07222__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_271_clk_i clknet_5_13__leaf_clk_i clknet_leaf_271_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_80_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_190_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08345_ _03967_ _01404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_80_83 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10784__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13160__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10284__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_173_3698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08276_ _03754_ memory\[18\]\[1\] _03929_ _03931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08254__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11679__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08229__I0 _03775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07227_ _03345_ _00908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_171_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_134_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11608__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_286_clk_i clknet_5_14__leaf_clk_i clknet_leaf_286_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_116_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10036__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07158_ _03298_ _00886_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_0_clk_i clknet_5_4__leaf_clk_i clknet_leaf_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07089_ _03260_ _00855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12504__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1061 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12489__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_22_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10024__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_224_clk_i clknet_5_27__leaf_clk_i clknet_leaf_224_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_83_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12810_ _05677_ _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13533__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13790_ _00829_ clknet_leaf_349_clk_i memory\[16\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_9_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12741_ memory\[40\]\[17\] memory\[41\]\[17\] memory\[42\]\[17\] memory\[43\]\[17\]
+ _06875_ _06326_ _02142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_4
XANTENNA__12661__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_800 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15460_ _00419_ clknet_leaf_316_clk_i memory\[53\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12672_ _06871_ _06872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_239_clk_i clknet_5_15__leaf_clk_i clknet_leaf_239_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14411_ _01450_ clknet_leaf_191_clk_i memory\[20\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12973__I _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08468__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11623_ memory\[32\]\[1\] memory\[33\]\[1\] memory\[34\]\[1\] memory\[35\]\[1\] _05742_
+ _05743_ _05838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15391_ _00350_ clknet_leaf_348_clk_i memory\[51\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_33_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06891__A2 _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14342_ _01381_ clknet_leaf_195_clk_i memory\[18\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06971__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_13_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_1323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11554_ memory\[28\]\[0\] memory\[29\]\[0\] _05769_ _05770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07140__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10505_ _05029_ memory\[4\]\[11\] _05156_ _05158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14273_ _01312_ clknet_leaf_414_clk_i memory\[29\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11485_ _03120_ _05701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_123_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09968__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13224_ _02213_ _02617_ _02352_ _02618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_33_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10436_ _05121_ _00261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_100_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_33_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_94_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07443__I1 _03336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13155_ memory\[32\]\[23\] memory\[33\]\[23\] memory\[34\]\[23\] memory\[35\]\[23\]
+ _02205_ _02345_ _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_10367_ _05026_ memory\[47\]\[10\] _05084_ _05085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12106_ _05669_ _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13086_ memory\[32\]\[22\] memory\[33\]\[22\] memory\[34\]\[22\] memory\[35\]\[22\]
+ _02205_ _02345_ _02482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
X_10298_ _03177_ _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_40_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12037_ _05732_ _06241_ _06243_ _06245_ _06246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_139_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10869__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13245__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13988_ _01027_ clknet_leaf_318_clk_i memory\[59\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_610 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15727_ _00686_ clknet_leaf_254_clk_i memory\[61\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12939_ _05653_ _02337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15658_ _00617_ clknet_leaf_255_clk_i memory\[5\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_138_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_138_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14609_ _01648_ clknet_leaf_95_clk_i memory\[26\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06882__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15589_ _00548_ clknet_leaf_319_clk_i memory\[57\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_172_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_185_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07977__I _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08130_ _03814_ memory\[15\]\[30\] _03818_ _03852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_16_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_161_819 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06881__I _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08074__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12955__A2 _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_860 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_4_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_79_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11499__I _05675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08061_ _03814_ memory\[12\]\[30\] _03751_ _03815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07012_ _03214_ _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10018__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12832__B _06482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_777 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07434__I1 _03327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07418__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08963_ _04227_ memory\[27\]\[21\] _04308_ _04310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07914_ _03153_ memory\[19\]\[9\] _03711_ _03721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08894_ _04273_ _01647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09633__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07845_ _03684_ _01187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12891__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07776_ _03150_ memory\[6\]\[8\] _03639_ _03648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07153__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09515_ _03177_ _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_155_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12994__S _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12643__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_175_3738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08048__I _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09446_ _04565_ _01907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_175_3749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_13_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_192_933 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_121_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12793__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09377_ _04233_ memory\[33\]\[24\] _04524_ _04529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08328_ _03806_ memory\[18\]\[26\] _03951_ _03958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_10_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07122__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08259_ _03921_ _01364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10009__I0 _04610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08712__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11270_ _05563_ _00653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_162_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_104_Left_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10221_ _04992_ _00175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07328__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10152_ _04616_ memory\[44\]\[20\] _04955_ _04956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11921__A3 _06116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10083_ _04896_ _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14960_ _01999_ clknet_leaf_71_clk_i memory\[37\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_163_clk_i clknet_5_28__leaf_clk_i clknet_leaf_163_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_46_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13911_ _00950_ clknet_leaf_135_clk_i memory\[11\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_96_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10689__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14891_ _01930_ clknet_leaf_52_clk_i memory\[35\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06936__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13842_ _00881_ clknet_leaf_117_clk_i memory\[13\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06966__I net16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08159__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07063__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13773_ _00812_ clknet_leaf_199_clk_i memory\[14\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_178_clk_i clknet_5_28__leaf_clk_i clknet_leaf_178_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_134_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08689__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10985_ _05031_ memory\[56\]\[12\] _05410_ _05413_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10496__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15512_ _00471_ clknet_leaf_384_clk_i memory\[54\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12724_ memory\[14\]\[17\] memory\[15\]\[17\] _06302_ _02125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15443_ _00402_ clknet_leaf_262_clk_i memory\[52\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12655_ memory\[12\]\[16\] memory\[13\]\[16\] _06714_ _06855_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_183_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_101_clk_i clknet_5_21__leaf_clk_i clknet_leaf_101_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11313__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11606_ memory\[6\]\[1\] memory\[7\]\[1\] _05706_ _05821_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15374_ _00333_ clknet_leaf_258_clk_i memory\[50\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12586_ memory\[8\]\[15\] memory\[9\]\[15\] memory\[10\]\[15\] memory\[11\]\[15\]
+ _06582_ _06721_ _06787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__07113__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_96_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14325_ _01364_ clknet_leaf_115_clk_i memory\[17\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_20_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11537_ _05752_ _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08861__I0 _04193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_123_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_53_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14256_ _01295_ clknet_leaf_114_clk_i memory\[15\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_116_clk_i clknet_5_23__leaf_clk_i clknet_leaf_116_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11468_ _05683_ _05684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA_clkbuf_leaf_323_clk_i_I clknet_5_10__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13207_ _02600_ _02601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_74_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10419_ _05112_ _00253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07416__I1 _03303_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14187_ _01226_ clknet_leaf_194_clk_i memory\[19\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12144__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11399_ _05632_ _00713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10176__A2 _04787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_21_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10420__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13138_ memory\[6\]\[23\] memory\[7\]\[23\] _02322_ _02533_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_5_28__f_clk_i clknet_2_3_0_clk_i clknet_5_28__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13069_ _06848_ _02464_ _06707_ _02465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__09453__S _04560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_119_Right_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__06927__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07630_ _03135_ memory\[10\]\[3\] _03567_ _03571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_109_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_1179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07561_ _03135_ memory\[0\]\[3\] _03530_ _03534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_157_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09300_ _04465_ _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_17_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07492_ memory\[59\]\[3\] _03315_ _03493_ _03497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07352__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09231_ _04451_ _01806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09162_ _04222_ memory\[30\]\[19\] _04405_ _04415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_84_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_170_3646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08113_ _03843_ _01296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_170_3657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12118__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09093_ _04378_ _01741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08044_ _03803_ _01267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1248 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08532__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13658__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12562__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08604__I0 _03810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_80_clk_i clknet_5_17__leaf_clk_i clknet_leaf_80_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12989__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09995_ _04595_ memory\[42\]\[10\] _04872_ _04873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11893__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_82 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08946_ _04210_ memory\[27\]\[13\] _04297_ _04301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_32_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_129_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08877_ _04264_ _01639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11667__A2 _05873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_95_clk_i clknet_5_20__leaf_clk_i clknet_leaf_95_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_4_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07828_ _03111_ memory\[7\]\[0\] _03675_ _03676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10302__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_93_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07759_ _03638_ _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_6_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10478__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07099__A2 net76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12711__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10770_ _05298_ _00418_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_67_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07611__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_410 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_272_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09429_ _04556_ _01899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11133__S _05482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_136_145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12440_ _06159_ _06642_ _06018_ _06643_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_81_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_666 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12371_ memory\[0\]\[12\] memory\[1\]\[12\] memory\[2\]\[12\] memory\[3\]\[12\] _06020_
+ _06090_ _06575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_23_817 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10972__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_33_clk_i clknet_5_7__leaf_clk_i clknet_leaf_33_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_22_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_112_Left_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_23_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14110_ _01149_ clknet_leaf_309_clk_i memory\[6\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09538__S _04617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11322_ memory\[61\]\[10\] _03155_ _05591_ _05592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07271__A2 _03264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15090_ _00049_ clknet_leaf_13_clk_i memory\[41\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_132_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_105_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14041_ _01080_ clknet_leaf_54_clk_i memory\[0\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_91_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11253_ _03329_ memory\[60\]\[10\] _05554_ _05555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_28_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10204_ _04983_ _00167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10402__I0 _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_48_clk_i clknet_5_18__leaf_clk_i clknet_leaf_48_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_52_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11184_ _05506_ _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_98_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10135_ _04600_ memory\[44\]\[12\] _04944_ _04947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09273__S _04466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09020__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14943_ _01982_ clknet_leaf_437_clk_i memory\[37\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10066_ _04910_ _00102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12855__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_121_Left_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14874_ _01913_ clknet_leaf_5_clk_i memory\[34\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07582__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13825_ _00864_ clknet_leaf_280_clk_i memory\[13\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13523__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_67_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13756_ _00795_ clknet_leaf_278_clk_i memory\[14\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08617__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10968_ _05014_ memory\[56\]\[4\] _05399_ _05404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_70_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07521__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12707_ memory\[52\]\[17\] memory\[53\]\[17\] _06832_ _02108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13687_ _03073_ _00762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10899_ _05367_ _00478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15426_ _00385_ clknet_leaf_316_clk_i memory\[52\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12638_ _05689_ _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_143_616 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_130_Left_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_31_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_370 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15357_ _00316_ clknet_leaf_347_clk_i memory\[50\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12569_ _06146_ _06769_ _06287_ _06770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__11594__A1 _05668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14308_ _01347_ clknet_leaf_368_clk_i memory\[17\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08352__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15288_ _00247_ clknet_leaf_386_clk_i memory\[47\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12218__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_180_1031 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14239_ _01278_ clknet_leaf_372_clk_i memory\[15\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08800_ _03174_ _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10944__I1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09780_ memory\[3\]\[6\] _03143_ _04751_ _04758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06992_ _03199_ _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XPHY_EDGE_ROW_7_Right_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09183__S _04416_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08731_ _03800_ memory\[24\]\[23\] _04168_ _04172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11649__A2 _05833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11726__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12846__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11218__S _05529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08662_ _04135_ _01553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10122__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_1_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07573__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07613_ _03212_ memory\[0\]\[28\] _03552_ _03561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_124_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08593_ _04098_ _01521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_152_1133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_178_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07544_ memory\[59\]\[28\] _03367_ _03515_ _03524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_793 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07475_ _03486_ _01015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09214_ _04206_ memory\[31\]\[11\] _04441_ _04443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_668 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09078__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_569 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09145_ _04406_ _01765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10792__S _05301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12621__I1 net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09358__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08262__S _03915_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09076_ _04203_ memory\[2\]\[10\] _04369_ _04370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_20_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11680__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08027_ _03791_ memory\[12\]\[19\] _03773_ _03792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10591__I _05180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_102_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_219_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11888__A2 _06098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_1267 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_590 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09978_ _04579_ memory\[42\]\[2\] _04861_ _04864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08929_ _04193_ memory\[27\]\[5\] _04286_ _04292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12837__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10699__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10032__S _04883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11940_ _05693_ _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_19_1103 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11871_ memory\[48\]\[5\] memory\[49\]\[5\] memory\[50\]\[5\] memory\[51\]\[5\] _06010_
+ _05694_ _06082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_67_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_98_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_39_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13610_ _02498_ _02997_ _05665_ _02998_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10822_ _05325_ _05326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_184_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14590_ _01629_ clknet_leaf_415_clk_i memory\[26\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08437__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_922 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13541_ _05690_ _02929_ _02930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_138_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10753_ _03266_ _03451_ _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_149_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_45_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_45_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10871__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13014__A1 _06720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09069__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13472_ _02337_ _02857_ _02859_ _02861_ _02862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12448__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10684_ _05252_ _00378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_70_709 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15211_ _00170_ clknet_leaf_36_clk_i memory\[45\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12423_ _06625_ _06626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_168_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15142_ _00101_ clknet_leaf_22_clk_i memory\[43\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12354_ memory\[62\]\[12\] memory\[63\]\[12\] _06557_ _06558_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11305_ memory\[61\]\[2\] _03131_ _05580_ _05583_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15073_ _00032_ clknet_leaf_438_clk_i memory\[41\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12285_ _03122_ _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_10_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10207__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14024_ _01063_ clknet_leaf_247_clk_i memory\[0\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_103_1308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11236_ _03313_ memory\[60\]\[2\] _05543_ _05546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09241__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11167_ _05509_ _00604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12422__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10118_ _04583_ memory\[44\]\[4\] _04933_ _04938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_175_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12828__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11098_ _03311_ memory\[58\]\[1\] _05471_ _05473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_145_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_22 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11038__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10049_ _04901_ _00094_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_69_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14926_ _01965_ clknet_leaf_64_clk_i memory\[36\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07555__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11351__I1 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_106_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10877__S _05348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14857_ _01896_ clknet_leaf_46_clk_i memory\[34\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_141_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_58_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_187_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_13808_ _00847_ clknet_leaf_116_clk_i memory\[16\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13253__A1 _02163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14788_ _01827_ clknet_leaf_397_clk_i memory\[32\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_102_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12377__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07251__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13739_ _03101_ _00786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_82_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13052__I _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_82_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13005__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07260_ memory\[39\]\[28\] _03367_ _03351_ _03368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10862__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_168_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07483__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07050__I _03228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_825 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07191_ _03143_ _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15409_ _00368_ clknet_leaf_156_clk_i memory\[51\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08807__I0 _04220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11501__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10614__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08082__S _03819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_1234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_123_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11300__I _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09901_ _04822_ _00025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_220_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09906__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08810__S _04204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10917__I1 _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_6_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09832_ memory\[3\]\[31\] _03220_ _04750_ _04785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_171_Right_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_165_3556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07426__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09763_ _04639_ memory\[38\]\[31\] _04713_ _04748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12819__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_06975_ _03186_ _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XTAP_TAPCELL_ROW_126_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08714_ _03783_ memory\[24\]\[15\] _04157_ _04163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_20_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09694_ _04711_ _02009_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07225__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09641__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08645_ _04126_ _01545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_90_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07171__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_516 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08576_ _04089_ _01513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13244__A1 _02592_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_77_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07161__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_37_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07527_ _03492_ _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_49_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07458_ memory\[49\]\[20\] _03350_ _03477_ _03478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_146_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_174_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07389_ _03439_ _00976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_150_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11411__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07895__I _03710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09088__S _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09128_ _04397_ _01757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_40_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_115_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_121_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09059_ _04187_ memory\[2\]\[2\] _04358_ _04361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09816__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12070_ _06276_ _06277_ _06001_ _06278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__08720__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10908__I1 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11030__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11021_ _05431_ _00536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09774__I1 _03134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_21_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12242__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output60_I net60 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07785__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07336__S _03401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15760_ _00719_ clknet_leaf_163_clk_i memory\[62\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12972_ _02369_ _02370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_86_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_86_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_422_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14711_ _01750_ clknet_leaf_58_clk_i memory\[2\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11923_ _06133_ _00736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10697__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15691_ _00650_ clknet_leaf_229_clk_i memory\[60\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13073__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_169_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_47_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_86_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14642_ _01681_ clknet_leaf_81_clk_i memory\[27\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13235__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11854_ _05794_ _06065_ _06066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__06974__I net19 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08167__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12197__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_64_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10805_ _05056_ memory\[53\]\[24\] _05312_ _05317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14573_ _01612_ clknet_leaf_125_clk_i memory\[25\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12589__A3 _06789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11785_ _05997_ _00734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11797__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13524_ _05772_ _02912_ _05775_ _02913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10844__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10736_ _05280_ _00402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_24_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13455_ memory\[0\]\[28\] memory\[1\]\[28\] memory\[2\]\[28\] memory\[3\]\[28\] _05784_
+ _03226_ _02845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10667_ memory\[51\]\[23\] _03196_ _05240_ _05244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11549__A1 _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13094__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12406_ _05667_ _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_35_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_619 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13386_ _05715_ _02772_ _02774_ _02776_ _02777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_106_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10598_ _05054_ memory\[50\]\[23\] _05203_ _05207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15125_ _00084_ clknet_leaf_10_clk_i memory\[42\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12337_ memory\[24\]\[11\] memory\[25\]\[11\] memory\[26\]\[11\] memory\[27\]\[11\]
+ _06472_ _05922_ _06542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_181_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09726__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15056_ _00015_ clknet_leaf_8_clk_i memory\[40\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09214__I0 _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12268_ _05921_ _06473_ _06474_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14007_ _01046_ clknet_leaf_261_clk_i memory\[59\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11219_ _05536_ _00629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12199_ _05794_ _06405_ _06406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_43_1295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07776__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09525__I _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_143_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_143_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_94_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_39_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_160_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__11324__I1 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13491__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14909_ _01948_ clknet_leaf_436_clk_i memory\[36\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_121_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08430_ _04000_ _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_77_127 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06884__I net2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10400__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_685 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13226__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_114_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_88 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_74_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11088__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08361_ _03975_ _01412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13321__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13711__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07312_ _03398_ _00940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10835__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_22_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08292_ _03770_ memory\[18\]\[9\] _03929_ _03939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07700__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07243_ _03356_ _00913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12327__S _05907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_969 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_119_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07174_ memory\[39\]\[0\] _03303_ _03309_ _03310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09453__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_160_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_44_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_371_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_184_3921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09205__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__S _04036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_371 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13158__S _02210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11012__I0 _05058_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12062__S _05802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_180_3829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09815_ _04776_ _02065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09746_ _04739_ _02033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06958_ net14 _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13465__A1 _02319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11315__I1 _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09371__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09677_ _04621_ memory\[37\]\[22\] _04700_ _04703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06889_ _03120_ _03121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__08192__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11406__S _05627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08628_ _04117_ _01537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08559_ _04080_ _01505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_37_514 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11205__I _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_42_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11570_ memory\[20\]\[0\] memory\[21\]\[0\] _05785_ _05786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10521_ _05045_ memory\[4\]\[19\] _05156_ _05166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_123_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_254 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_468 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13240_ memory\[16\]\[24\] memory\[17\]\[24\] memory\[18\]\[24\] memory\[19\]\[24\]
+ _02233_ _02376_ _02634_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_17_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_91_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10452_ _05129_ _00269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_116_991 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13171_ _02501_ _02565_ _02566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10383_ _05043_ memory\[47\]\[18\] _05084_ _05093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11951__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12122_ _05731_ _06317_ _06329_ _06330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_102_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13068__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12053_ memory\[20\]\[7\] memory\[21\]\[7\] _05785_ _06262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_116_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11004_ _05050_ memory\[56\]\[21\] _05421_ _05423_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15812_ _00771_ clknet_leaf_299_clk_i memory\[9\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12700__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13456__A1 _05759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15743_ _00702_ clknet_leaf_310_clk_i memory\[62\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12955_ _02213_ _02351_ _02352_ _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_29_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_59_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_29_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11906_ memory\[28\]\[5\] memory\[29\]\[5\] _05915_ _06117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_1255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_1266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10220__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12886_ memory\[28\]\[19\] memory\[29\]\[19\] _06604_ _02285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15674_ _00633_ clknet_leaf_396_clk_i memory\[5\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13303__S1 _02376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14625_ _01664_ clknet_leaf_416_clk_i memory\[27\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11837_ memory\[40\]\[4\] memory\[41\]\[4\] memory\[42\]\[4\] memory\[43\]\[4\] _05761_
+ _05762_ _06049_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
Xclkbuf_leaf_407_clk_i clknet_5_3__leaf_clk_i clknet_leaf_407_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_7_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13531__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_322 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10817__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14556_ _01595_ clknet_leaf_390_clk_i memory\[25\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_138_571 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11768_ memory\[28\]\[3\] memory\[29\]\[3\] _05915_ _05981_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08625__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09683__I0 _04627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13507_ _02895_ _02896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10719_ _05271_ _00394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14487_ _01526_ clknet_leaf_105_clk_i memory\[22\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_70_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11699_ _05731_ _05904_ _05912_ _05913_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__11051__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_3_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_13438_ memory\[62\]\[28\] memory\[63\]\[28\] _02448_ _02828_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_126_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_753 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_180_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_449 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11242__I0 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13369_ _02358_ _02753_ _02760_ _02761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_0_140_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11942__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_77_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15108_ _00067_ clknet_leaf_442_clk_i memory\[42\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08360__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07930_ _03729_ _01227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15039_ _02078_ clknet_leaf_439_clk_i memory\[40\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__06879__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_162_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12042__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07861_ _03175_ memory\[7\]\[16\] _03686_ _03693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_177_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__15382__CLK clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09600_ _04612_ memory\[36\]\[18\] _04653_ _04662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13706__S _03075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07792_ _03656_ _01162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_3_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_39_1139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07704__S _03603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09191__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09531_ _03193_ _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_155_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_155_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11226__S _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09462_ _03305_ _03376_ _04574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA_clkbuf_leaf_318_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_622 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07921__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_650 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08413_ _04003_ _01436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_148_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09393_ _03305_ net72 _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_177_3780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08344_ _03754_ memory\[1\]\[1\] _03965_ _03967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_62_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10864__I _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08275_ _03930_ _01371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_173_3699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07226_ memory\[39\]\[17\] _03344_ _03330_ _03345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09426__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11608__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12186__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07157_ _03209_ memory\[13\]\[27\] _03290_ _03298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_30_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09366__S _04513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08270__S _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07088_ _03212_ memory\[16\]\[28\] _03251_ _03260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11909__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10305__S _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_1211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13150__A3 _02544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13616__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11644__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09729_ _04730_ _02025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13533__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08165__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12740_ _06322_ _02140_ _06461_ _02141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_26_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_26_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07912__I0 _03150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12671_ memory\[44\]\[16\] memory\[45\]\[16\] _06319_ _06871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14410_ _01449_ clknet_leaf_192_clk_i memory\[20\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11622_ _05736_ _05836_ _05739_ _05837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_108_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15390_ _00349_ clknet_leaf_348_clk_i memory\[51\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_37_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08445__S _04012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13610__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_13_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14341_ _01380_ clknet_leaf_366_clk_i memory\[18\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_42_clk_i_I clknet_5_18__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11553_ _05655_ _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_108_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_393_clk_i clknet_5_6__leaf_clk_i clknet_leaf_393_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10504_ _05157_ _00293_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14272_ _01311_ clknet_leaf_354_clk_i memory\[29\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_98_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11484_ _05653_ _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_162_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12177__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13223_ memory\[46\]\[24\] memory\[47\]\[24\] _02487_ _02617_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11224__I0 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10435_ _05026_ memory\[48\]\[10\] _05120_ _05121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_59_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08180__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13154_ _02341_ _02548_ _06866_ _02549_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10366_ _05072_ _05084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08640__I1 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12105_ _05736_ _06312_ _06177_ _06313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_104_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10215__S _04980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13085_ _02341_ _02480_ _06866_ _02481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_10297_ _05040_ _00203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_267_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09075__I _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12036_ _05741_ _06244_ _06245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_72_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_40_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_331_clk_i clknet_5_10__leaf_clk_i clknet_leaf_331_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_176_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13987_ _01026_ clknet_leaf_321_clk_i memory\[59\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08156__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12101__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11046__S _05435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15726_ _00685_ clknet_leaf_255_clk_i memory\[61\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12938_ _03304_ _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_34_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_346_clk_i clknet_5_8__leaf_clk_i clknet_leaf_346_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_34_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_29_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_185_430 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15657_ _00616_ clknet_leaf_246_clk_i memory\[5\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10885__S _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12869_ _06713_ _02263_ _02265_ _02267_ _02268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_75_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13288__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_186_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_138_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14608_ _01647_ clknet_leaf_97_clk_i memory\[26\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09656__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15588_ _00547_ clknet_leaf_319_clk_i memory\[57\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14539_ _01578_ clknet_leaf_187_clk_i memory\[24\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_141_67 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_79_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_160_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_116_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08060_ _03217_ _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XTAP_TAPCELL_ROW_116_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_1080 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07011_ net28 _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__12605__S _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11729__B _05939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08631__I1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_266 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08962_ _04309_ _01679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13668__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09914__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07913_ _03720_ _01219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08893_ _04224_ memory\[26\]\[20\] _04272_ _04273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_16_Left_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_75_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07198__I1 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_62 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13436__S _05702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12340__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07844_ _03150_ memory\[7\]\[8\] _03675_ _03684_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07434__S _03455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07775_ _03647_ _01154_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_179_3820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09514_ _04609_ _01931_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12643__A2 _06830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_91_1174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09445_ _04233_ memory\[34\]\[24\] _04560_ _04565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_52_1147 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_175_3739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_137_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09376_ _04528_ _01874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_191_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09647__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08327_ _03957_ _01396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_10_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_7_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_488 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08258_ _03804_ memory\[17\]\[25\] _03915_ _03921_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_127_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_160_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11206__I0 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07209_ _03333_ _00902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_166_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08189_ _03884_ _01331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_43_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07609__S _03552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10220_ _04616_ memory\[45\]\[20\] _04991_ _04992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_123_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_37_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10151_ _04932_ _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_30_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11921__A4 _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_63_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13203__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09824__S _04773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10082_ _04918_ _00110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08386__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07189__I1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12331__A1 _06318_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13910_ _00949_ clknet_leaf_134_clk_i memory\[11\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14890_ _01929_ clknet_leaf_45_clk_i memory\[35\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_50_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07344__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13841_ _00880_ clknet_leaf_118_clk_i memory\[13\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08138__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13772_ _00811_ clknet_leaf_199_clk_i memory\[14\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09886__I0 _04623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10984_ _05412_ _00518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_69_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15511_ _00470_ clknet_leaf_383_clk_i memory\[54\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12723_ _02123_ _02124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12984__I _03122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12654_ _06844_ _06847_ _06850_ _06853_ _06854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15442_ _00401_ clknet_leaf_263_clk_i memory\[52\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08175__S _03868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13434__I1 net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12398__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11605_ _05819_ _05820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_167_1024 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12585_ _06717_ _06785_ _06304_ _06786_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12937__A3 _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_174 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08066__A2 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15373_ _00332_ clknet_leaf_257_clk_i memory\[50\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14324_ _01363_ clknet_leaf_104_clk_i memory\[17\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11536_ _03118_ _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08903__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12933__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_151_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_68_1176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14255_ _01294_ clknet_leaf_171_clk_i memory\[15\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11467_ _03119_ _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XTAP_TAPCELL_ROW_150_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_123_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_886 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13206_ memory\[12\]\[24\] memory\[13\]\[24\] _05769_ _02600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07519__S _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10418_ _05010_ memory\[48\]\[2\] _05109_ _05112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14186_ _01225_ clknet_leaf_207_clk_i memory\[19\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_21_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_74_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_396 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11398_ _03338_ memory\[62\]\[14\] _05627_ _05632_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_111_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13137_ _02531_ _02532_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_103_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10349_ _05075_ _00220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_104_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09734__S _04725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_270_clk_i clknet_5_13__leaf_clk_i clknet_leaf_270_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13068_ memory\[6\]\[22\] memory\[7\]\[22\] _02322_ _02464_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08377__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13256__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12019_ _06159_ _06227_ _06018_ _06228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_174_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10184__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07254__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_285_clk_i clknet_5_14__leaf_clk_i clknet_leaf_285_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07560_ _03533_ _01053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09877__I0 _04614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_157_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15709_ _00668_ clknet_leaf_336_clk_i memory\[61\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_75_203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07491_ _03496_ _01021_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_158_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09230_ _04222_ memory\[31\]\[19\] _04441_ _04451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_158_485 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_115_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_173_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09161_ _04414_ _01773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_146_669 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08301__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13681__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08112_ _03796_ memory\[15\]\[21\] _03841_ _03843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_170_3647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09092_ _04220_ memory\[2\]\[18\] _04369_ _04378_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_32_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_475 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08043_ _03802_ memory\[12\]\[24\] _03794_ _03803_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_223_clk_i clknet_5_27__leaf_clk_i clknet_leaf_223_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_131_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12335__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12134__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09994_ _04860_ _04872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_50_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__07228__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_86_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_238_clk_i clknet_5_26__leaf_clk_i clknet_leaf_238_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_86_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_110_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08945_ _04300_ _01671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12313__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13166__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_23_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_32_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08876_ _04208_ memory\[26\]\[12\] _04261_ _04264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_input22_I data_i[23] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07040__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07827_ _03674_ _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_98_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_717 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_93_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07758_ _03124_ _03528_ _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_79_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_79_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07689_ _03601_ _01114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_215_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08540__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_66_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09428_ _04216_ memory\[34\]\[16\] _04549_ _04556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11427__I0 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09359_ _04519_ _01866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_81_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_180_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_152_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12370_ _06159_ _06573_ _06018_ _06574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_63_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_133_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_829 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_185_Right_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_34_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11321_ _05579_ _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_133_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12245__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10650__I1 _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14040_ _01079_ clknet_leaf_55_clk_i memory\[0\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11252_ _05542_ _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_91_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_24_1013 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10203_ _04600_ memory\[45\]\[12\] _04980_ _04983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_11183_ _05517_ _00612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_52_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10134_ _04946_ _00134_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_1079 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_41_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14942_ _01981_ clknet_leaf_435_clk_i memory\[37\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10065_ _04598_ memory\[43\]\[11\] _04908_ _04910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10166__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07074__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14873_ _01912_ clknet_leaf_70_clk_i memory\[34\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13824_ _00863_ clknet_leaf_279_clk_i memory\[13\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09859__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07802__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10967_ _05403_ _00510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13755_ _03109_ _00794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07334__I1 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11324__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11910__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_104_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12706_ _06272_ _02102_ _02104_ _02106_ _02107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_155_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10898_ memory\[55\]\[3\] _03134_ _05363_ _05367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13686_ _03072_ net64 _03122_ _03073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_39_984 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15425_ _00384_ clknet_leaf_329_clk_i memory\[52\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12637_ _06835_ _06836_ _06287_ _06837_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_38_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15356_ _00315_ clknet_leaf_346_clk_i memory\[50\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08633__S _04110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12568_ memory\[54\]\[15\] memory\[55\]\[15\] _06421_ _06769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_0_1162 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_2_1_0_clk_i clknet_0_clk_i clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_152_Right_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14307_ _01346_ clknet_leaf_342_clk_i memory\[17\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11519_ _05734_ _05735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_13_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15287_ _00246_ clknet_leaf_39_clk_i memory\[47\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12218__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12499_ _06149_ _06700_ _06701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_417_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09528__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14238_ _01277_ clknet_leaf_372_clk_i memory\[15\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_536 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08598__I0 _03804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12543__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_145_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11977__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14169_ _01208_ clknet_leaf_54_clk_i memory\[7\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_1184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__09464__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06991_ net23 _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_164_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08730_ _04171_ _01585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__06887__I net1 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11649__A3 _05848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08661_ memory\[23\]\[22\] _03355_ _04132_ _04135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07612_ _03560_ _01078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08770__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08592_ _03798_ memory\[22\]\[22\] _04095_ _04098_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_156_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_124_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_63 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07543_ _03523_ _01046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08522__I0 _03796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11234__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07474_ memory\[49\]\[28\] _03367_ _03477_ _03486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_118_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_48_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09213_ _04442_ _01797_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_88_1316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_107_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_134_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09144_ _04203_ memory\[30\]\[10\] _04405_ _04406_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_162_clk_i clknet_5_25__leaf_clk_i clknet_leaf_162_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_17_656 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09639__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_98_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA_clkbuf_leaf_89_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_138 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11585__A2 _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_16_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_71_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12782__A1 _06831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09075_ _04357_ _04369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_142_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_875 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07159__S _03290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08026_ _03183_ _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_47_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_187_3963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_177_clk_i clknet_5_28__leaf_clk_i clknet_leaf_177_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12385__I1 memory\[39\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_60_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10396__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09977_ _04863_ _00060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_100_clk_i clknet_5_21__leaf_clk_i clknet_leaf_100_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08928_ _04291_ _01663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12837__A2 _02228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07013__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08859_ _04191_ memory\[26\]\[4\] _04250_ _04255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08761__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11870_ _05682_ _06080_ _05687_ _06081_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_54_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08718__S _04157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12748__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_115_clk_i clknet_5_23__leaf_clk_i clknet_leaf_115_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10821_ _03124_ _03451_ _05325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08513__I0 _03787_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11144__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_366_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10752_ _05288_ _00410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13540_ memory\[40\]\[29\] memory\[41\]\[29\] memory\[42\]\[29\] memory\[43\]\[29\]
+ _05692_ _05694_ _02929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_39_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_95_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_95_898 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_45_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_45_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_397 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13471_ _02344_ _02860_ _02861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_164_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09069__I1 memory\[2\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10683_ memory\[51\]\[31\] _03220_ _05217_ _05252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_82_548 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10983__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12448__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15210_ _00169_ clknet_leaf_38_clk_i memory\[45\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12422_ memory\[60\]\[13\] memory\[61\]\[13\] _06273_ _06625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_62_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12773__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12353_ _05661_ _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10623__I1 _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15141_ _00100_ clknet_leaf_445_clk_i memory\[43\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_121_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07069__S _03240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_161_992 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11304_ _05582_ _00668_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_51_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15072_ _00031_ clknet_leaf_437_clk_i memory\[41\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12284_ _06427_ _06444_ _06466_ _06489_ _06490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_14023_ _01062_ clknet_leaf_246_clk_i memory\[0\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11235_ _05545_ _00636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09284__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11166_ _03311_ memory\[5\]\[1\] _05507_ _05509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11319__S _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10117_ _04937_ _00126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11097_ _05472_ _00571_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10139__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10048_ _04581_ memory\[43\]\[3\] _04897_ _04901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14925_ _01964_ clknet_leaf_49_clk_i memory\[36\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_69_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08752__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_300 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14856_ _01895_ clknet_leaf_45_clk_i memory\[34\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_193_4112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_141_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12658__B _06304_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07532__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13807_ _00846_ clknet_leaf_194_clk_i memory\[16\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_14787_ _01826_ clknet_leaf_403_clk_i memory\[32\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_534 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07307__I1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11999_ _06208_ net68 _05802_ _06209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13738_ _03357_ memory\[9\]\[23\] _03097_ _03101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_82_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_128_433 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13005__A2 _02401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13669_ _03304_ _03048_ _03055_ _03056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_128_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13636__S0 _05725_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_183_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_13_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09459__S _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15408_ _00367_ clknet_leaf_153_clk_i memory\[51\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08363__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07190_ _03320_ _00896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_155_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_90_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_5_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_87_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15339_ _00298_ clknet_leaf_244_clk_i memory\[4\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_94_clk_i clknet_5_20__leaf_clk_i clknet_leaf_94_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_13_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09258__I _04465_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09900_ _04637_ memory\[40\]\[30\] _04788_ _04822_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_111_377 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_10_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_165_3546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09831_ _04784_ _02073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_165_3557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08991__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_5_12__f_clk_i clknet_2_1_0_clk_i clknet_5_12__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10133__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09762_ _04747_ _02041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06974_ net19 _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_182_3882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_20_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07506__I _03492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09922__S _04825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_119_1305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08713_ _04162_ _01577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09693_ _04637_ memory\[37\]\[30\] _04677_ _04711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_32_clk_i clknet_5_7__leaf_clk_i clknet_leaf_32_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08743__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__I1 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08644_ memory\[23\]\[14\] _03338_ _04121_ _04126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08538__S _04059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10550__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__12127__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07171__A2 _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11472__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08575_ _03781_ memory\[22\]\[14\] _04084_ _04089_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13244__A2 _02607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07526_ _03514_ _01038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10302__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_47_clk_i clknet_5_18__leaf_clk_i clknet_leaf_47_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_119_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07241__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_932 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07457_ _03454_ _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_18_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09369__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_902 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07388_ _03191_ memory\[8\]\[21\] _03437_ _03439_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_134_436 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12755__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_17_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09127_ _04187_ memory\[30\]\[2\] _04394_ _04397_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_161_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_40_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09058_ _04360_ _01724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_102_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_642 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_856 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08009_ _03779_ memory\[12\]\[13\] _03773_ _03780_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_8_Left_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__10369__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13180__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_1077 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07617__S _03529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11020_ _05066_ memory\[56\]\[29\] _05421_ _05431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08800__I _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_25_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output53_I net53 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09832__S _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12971_ memory\[20\]\[20\] memory\[21\]\[20\] _02368_ _02369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10978__S _05399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14710_ _01749_ clknet_leaf_59_clk_i memory\[2\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_86_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11922_ _06132_ net67 _05802_ _06133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15690_ _00649_ clknet_leaf_229_clk_i memory\[60\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07352__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_47_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14641_ _01680_ clknet_leaf_95_clk_i memory\[27\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11853_ memory\[16\]\[4\] memory\[17\]\[4\] memory\[18\]\[4\] memory\[19\]\[4\] _05795_
+ _05796_ _06065_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_86_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_848 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10804_ _05316_ _00434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14572_ _01611_ clknet_leaf_186_clk_i memory\[25\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08247__I _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11784_ _05996_ net65 _05802_ _05997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_112_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13523_ memory\[14\]\[29\] memory\[15\]\[29\] _05773_ _02912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10735_ _05054_ memory\[52\]\[23\] _05276_ _05280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_24_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13618__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_153_723 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_82_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13454_ _05752_ _02843_ _05791_ _02844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_70_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10666_ _05243_ _00369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_24_924 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13094__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12405_ _06607_ _06608_ _06195_ _06609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_153_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13385_ _05724_ _02775_ _02776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10597_ _05206_ _00337_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_24_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_765 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15124_ _00083_ clknet_leaf_10_clk_i memory\[42\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12336_ _05918_ _06540_ _06195_ _06541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__08911__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12349__I1 net42 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13529__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12267_ memory\[24\]\[10\] memory\[25\]\[10\] memory\[26\]\[10\] memory\[27\]\[10\]
+ _06472_ _05922_ _06473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_50_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15055_ _00014_ clknet_leaf_19_clk_i memory\[40\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_103_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13171__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_697 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14006_ _01045_ clknet_leaf_160_clk_i memory\[59\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11218_ _03363_ memory\[5\]\[26\] _05529_ _05536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12198_ memory\[16\]\[9\] memory\[17\]\[9\] memory\[18\]\[9\] memory\[19\]\[9\] _06342_
+ _05796_ _06405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__11049__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08973__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11149_ _05499_ _00596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_143_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_1337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10780__I0 _05031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_37_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_160_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08725__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07528__I1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13264__S _02322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14908_ _01947_ clknet_leaf_435_clk_i memory\[36\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10532__I0 _05056_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08358__S _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_156_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_144_45 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_176_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_506 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14839_ _01878_ clknet_leaf_73_clk_i memory\[33\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08360_ _03770_ memory\[1\]\[9\] _03965_ _03975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_15_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_07311_ memory\[11\]\[17\] _03344_ _03390_ _03398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09150__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08291_ _03938_ _01379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_73_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07242_ memory\[39\]\[22\] _03355_ _03351_ _03356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08093__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1000 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_6_645 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_119_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13012__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12407__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07173_ _03308_ _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_119_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10128__S _04933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12851__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_314_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_184_3911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_111_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_10_651 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07437__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09814_ memory\[3\]\[22\] _03193_ _04773_ _04776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_22_1358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10771__I0 _05022_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09652__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09745_ _04621_ memory\[38\]\[22\] _04736_ _04739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06957_ _03173_ _00810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07519__I1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08716__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08268__S _03892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09676_ _04702_ _02000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_97_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06888_ _03119_ _03120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_69_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_90_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12298__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08627_ memory\[23\]\[6\] _03321_ _04110_ _04117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08067__I _03818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08558_ _03764_ memory\[22\]\[6\] _04073_ _04080_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07900__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09141__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12976__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12520__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07509_ memory\[59\]\[11\] _03332_ _03504_ _03506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08489_ _04043_ _01472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_42_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09099__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10520_ _05165_ _00301_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_91_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_211 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_52_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12728__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_99_Left_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10451_ _05043_ memory\[48\]\[18\] _05120_ _05129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10038__S _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_150_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13170_ memory\[24\]\[23\] memory\[25\]\[23\] memory\[26\]\[23\] memory\[27\]\[23\]
+ _02363_ _02502_ _02565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08731__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10382_ _05092_ _00236_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12121_ _06318_ _06321_ _06324_ _06328_ _06329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__13349__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12052_ _05914_ _06256_ _06258_ _06260_ _06261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_2_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_57_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12900__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11003_ _05422_ _00527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_15811_ _00770_ clknet_leaf_302_clk_i memory\[9\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13084__S _06728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1235 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13700__I0 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15742_ _00701_ clknet_leaf_310_clk_i memory\[62\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_137_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12954_ _05664_ _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__07082__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_29_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11905_ _05731_ _06108_ _06115_ _06116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_59_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15673_ _00632_ clknet_leaf_152_clk_i memory\[5\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12885_ _06445_ _02276_ _02283_ _02284_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_14624_ _01663_ clknet_leaf_415_clk_i memory\[27\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_971 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11836_ _05753_ _06047_ _05757_ _06048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_114_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_150 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12967__A1 _06610_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07810__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_263_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14555_ _01594_ clknet_leaf_4_clk_i memory\[24\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_184_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11767_ _05731_ _05972_ _05979_ _05980_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_166_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11332__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13506_ memory\[52\]\[29\] memory\[53\]\[29\] _05716_ _02895_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07694__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10718_ _05037_ memory\[52\]\[15\] _05265_ _05271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14486_ _01525_ clknet_leaf_91_clk_i memory\[22\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11698_ _05748_ _05906_ _05909_ _05911_ _05912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_71_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13437_ _02826_ _02827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_113_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10649_ _05234_ _00361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_109_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13368_ _02367_ _02755_ _02757_ _02759_ _02760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_23_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15107_ _00066_ clknet_leaf_434_clk_i memory\[42\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_77_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12319_ _06523_ _06524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XTAP_TAPCELL_ROW_114_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13299_ memory\[20\]\[25\] memory\[21\]\[25\] _02368_ _02692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09199__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07257__S _03351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_139_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_15038_ _02077_ clknet_leaf_440_clk_i memory\[40\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_162_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08946__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07860_ _03692_ _01194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_78_1123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07791_ _03172_ memory\[6\]\[15\] _03650_ _03656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_20 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_78_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11458__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09530_ _04620_ _01936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__10505__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09371__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09461_ _03110_ _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_91_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08412_ _03754_ memory\[20\]\[1\] _04001_ _04003_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_114_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09392_ _04536_ _01882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_87_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09123__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12958__A1 _02209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_148_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08343_ _03966_ _01403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_175_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11242__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_879 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08274_ _03746_ memory\[18\]\[0\] _03929_ _03930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07225_ _03177_ _03344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_105_918 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_104_417 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_61 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09647__S _04678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13383__A1 _05719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07156_ _03297_ _00885_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11976__I _05691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07087_ _03259_ _00854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_112_461 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_100_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13135__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08937__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11697__A1 _05760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12801__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_29_Right_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_07989_ _03146_ _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__11417__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10321__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09728_ _04604_ memory\[38\]\[14\] _04725_ _04730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09362__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_409 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12741__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_26_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09659_ _04693_ _01992_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13632__S _05716_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_171_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12670_ _06446_ _06864_ _06867_ _06869_ _06870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_33_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07630__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11621_ memory\[38\]\[1\] memory\[39\]\[1\] _05737_ _05836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_77_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11152__S _05493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07676__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14340_ _01379_ clknet_leaf_367_clk_i memory\[18\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_181_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11552_ _05675_ _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_135_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_38_Right_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_162_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10503_ _05026_ memory\[4\]\[10\] _05156_ _05157_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14271_ _01310_ clknet_leaf_351_clk_i memory\[29\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11483_ _03114_ _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_98_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10991__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13222_ _02615_ _02616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10434_ _05108_ _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_59_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13587__B _05775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10365_ _05083_ _00228_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13153_ memory\[38\]\[23\] memory\[39\]\[23\] _06728_ _02548_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_143_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_21_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10983__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13126__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12104_ memory\[38\]\[8\] memory\[39\]\[8\] _06039_ _06312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13084_ memory\[38\]\[22\] memory\[39\]\[22\] _06728_ _02480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10296_ _05039_ memory\[46\]\[16\] _05027_ _05040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12035_ memory\[32\]\[7\] memory\[33\]\[7\] memory\[34\]\[7\] memory\[35\]\[7\] _05742_
+ _05743_ _06244_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_72_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10735__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_47_Right_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09292__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13986_ _01025_ clknet_leaf_320_clk_i memory\[59\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_87_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15725_ _00684_ clknet_leaf_244_clk_i memory\[61\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_158_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12937_ _02319_ _02327_ _02334_ _02335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_34_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_0_clk_i_I clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11160__I0 _03373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_87_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_150_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_407 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15656_ _00615_ clknet_leaf_245_clk_i memory\[5\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_34_1037 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12868_ _06720_ _02266_ _02267_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_157_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_146_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09105__I0 _04233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13288__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07540__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14607_ _01646_ clknet_leaf_124_clk_i memory\[26\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_138_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11819_ _05689_ _06031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_29_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15587_ _00546_ clknet_leaf_321_clk_i memory\[57\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_7_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12799_ _06713_ _02192_ _02196_ _02198_ _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XPHY_EDGE_ROW_56_Right_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_7_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_157_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14538_ _01577_ clknet_leaf_187_clk_i memory\[24\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_155_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_44_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_391 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_71_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_79_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14469_ _01508_ clknet_leaf_364_clk_i memory\[22\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_116_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07010_ _03213_ _00823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_126_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13365__A1 _02371_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09467__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08371__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_113_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_269 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_1193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10406__S _05095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10974__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13117__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08961_ _04224_ memory\[27\]\[20\] _04308_ _04309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_11_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08919__I0 _04181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_65_Right_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13717__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07912_ _03150_ memory\[19\]\[8\] _03711_ _03720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12621__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08892_ _04249_ _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10726__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08544__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07715__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09592__I0 _04604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07843_ _03683_ _01186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_79_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10141__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07774_ _03147_ memory\[6\]\[7\] _03639_ _03647_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_179_3810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09513_ _04608_ memory\[35\]\[16\] _04596_ _04609_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_908 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09444_ _04564_ _01906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_66_418 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08546__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_166_Right_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_EDGE_ROW_74_Right_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_192_913 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09375_ _04231_ memory\[33\]\[23\] _04524_ _04528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_46_131 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_434 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_6_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08326_ _03804_ memory\[18\]\[25\] _03951_ _03957_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11603__A1 _05651_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_159_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_10_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_34_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08257_ _03920_ _01363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_7_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_144_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_90_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_540 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07208_ memory\[39\]\[11\] _03332_ _03330_ _03333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09377__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08188_ _03802_ memory\[29\]\[24\] _03879_ _03884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07139_ _03288_ _00877_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_37_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13108__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_5_9__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_83_Right_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_93_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10150_ _04954_ _00142_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_211_clk_i_I clknet_5_27__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07830__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13203__S1 _06779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_406_clk_i clknet_5_3__leaf_clk_i clknet_leaf_406_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13627__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10081_ _04614_ memory\[43\]\[19\] _04908_ _04918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11390__I0 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_50_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13840_ _00879_ clknet_leaf_120_clk_i memory\[13\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09335__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_718 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09840__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13771_ _00810_ clknet_leaf_201_clk_i memory\[14\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_134_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11142__I0 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10983_ _05029_ memory\[56\]\[11\] _05410_ _05412_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13362__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15510_ _00469_ clknet_leaf_41_clk_i memory\[54\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_92_Right_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12722_ memory\[12\]\[17\] memory\[13\]\[17\] _06714_ _02123_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_139_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08456__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07360__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_133_Right_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15441_ _00400_ clknet_leaf_261_clk_i memory\[52\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12653_ _06851_ _06852_ _06853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_38_643 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_946 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_423 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07649__I0 _03163_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13595__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11604_ memory\[4\]\[1\] memory\[5\]\[1\] _05702_ _05819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_1092 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15372_ _00331_ clknet_leaf_272_clk_i memory\[50\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12584_ memory\[14\]\[15\] memory\[15\]\[15\] _06302_ _06785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_52_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_25_326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14323_ _01362_ clknet_leaf_102_clk_i memory\[17\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_128_1009 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11535_ _05750_ _05751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_68_1144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_184_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14254_ _01293_ clknet_leaf_197_clk_i memory\[15\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11466_ _05681_ _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_150_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_145_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13205_ _06844_ _02594_ _02596_ _02598_ _02599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__12505__I _05686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10417_ _05111_ _00252_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08074__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_74_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14185_ _01224_ clknet_leaf_206_clk_i memory\[19\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11397_ _05631_ _00712_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_74_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10226__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09810__I1 _03186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13136_ memory\[4\]\[23\] memory\[5\]\[23\] _06845_ _02531_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10348_ _05008_ memory\[47\]\[1\] _05073_ _05075_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13067_ _02462_ _02463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_10279_ _05028_ _00197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10708__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12018_ memory\[6\]\[7\] memory\[7\]\[7\] _05706_ _06227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11381__I0 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11057__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12240__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_178_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_109_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_109_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_413_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10896__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13969_ _01008_ clknet_leaf_158_clk_i memory\[49\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11133__I0 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15708_ _00667_ clknet_leaf_335_clk_i memory\[61\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07888__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07490_ memory\[59\]\[2\] _03313_ _03493_ _03496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_453 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_111_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_100_Right_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_15639_ _00598_ clknet_leaf_158_clk_i memory\[58\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_174_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09160_ _04220_ memory\[30\]\[18\] _04405_ _04414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_150_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_160_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_613 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_111_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_467 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08111_ _03842_ _01295_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13681__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_161_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09091_ _04377_ _01740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13338__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08042_ _03199_ _03802_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09197__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_47_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_131_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_4_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_589 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13020__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09801__I1 _03174_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07812__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09993_ _04871_ _00068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_110_784 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08944_ _04208_ memory\[27\]\[12\] _04297_ _04300_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12351__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09565__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07445__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_32_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08875_ _04263_ _01638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_99_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_1204 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_85_clk_i_I clknet_5_17__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_392_clk_i clknet_5_3__leaf_clk_i clknet_leaf_392_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07826_ _03306_ _03528_ _03674_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_93_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07244__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input15_I data_i[17] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09660__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09317__I0 _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07757_ _03637_ _01146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13182__S _02382_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11824__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08276__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07688_ _03221_ memory\[10\]\[31\] _03566_ _03601_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07180__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09427_ _04555_ _01898_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_137_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_19_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_165_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09358_ _04214_ memory\[33\]\[15\] _04513_ _04519_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_624 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08309_ _03787_ memory\[18\]\[17\] _03940_ _03948_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_330_clk_i clknet_5_10__leaf_clk_i clknet_leaf_330_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09289_ _04482_ _01833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_95_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11320_ _05590_ _00676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08803__I _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11251_ _05553_ _00644_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10046__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_30_340 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_91_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10202_ _04982_ _00166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_345_clk_i clknet_5_8__leaf_clk_i clknet_leaf_345_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_362_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11182_ _03327_ memory\[5\]\[9\] _05507_ _05517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_105_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13188__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13357__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10133_ _04598_ memory\[44\]\[11\] _04944_ _04946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_140_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__09556__I0 _04637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14941_ _01980_ clknet_leaf_435_clk_i memory\[37\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10064_ _04909_ _00101_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14872_ _01911_ clknet_leaf_69_clk_i memory\[34\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13823_ _00862_ clknet_leaf_373_clk_i memory\[13\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_3_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_35_Left_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13092__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08186__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13754_ _03373_ memory\[9\]\[31\] _03074_ _03109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10966_ _05012_ memory\[56\]\[3\] _05399_ _05403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07090__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_67_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_151_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_104_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12705_ _06279_ _02105_ _02106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_191_4040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11910__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_191_4051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13685_ _03026_ _03041_ _03056_ _03071_ _03072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_10897_ _05366_ _00477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15424_ _00383_ clknet_leaf_330_clk_i memory\[52\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13568__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_127_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12636_ memory\[54\]\[16\] memory\[55\]\[16\] _06421_ _06836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_122_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_152_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08295__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15355_ _00314_ clknet_leaf_392_clk_i memory\[4\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12567_ _06767_ _06768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_108_372 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11340__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14306_ _01345_ clknet_leaf_343_clk_i memory\[17\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09809__I _04750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11518_ memory\[36\]\[0\] memory\[37\]\[0\] _05733_ _05734_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15286_ _00245_ clknet_leaf_40_clk_i memory\[47\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12498_ memory\[48\]\[14\] memory\[49\]\[14\] memory\[50\]\[14\] memory\[51\]\[14\]
+ _06699_ _06150_ _06700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_1_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_44_Left_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14237_ _01276_ clknet_leaf_278_clk_i memory\[15\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11449_ _05664_ _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_46_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09745__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11977__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14168_ _01207_ clknet_leaf_53_clk_i memory\[7\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13119_ _02514_ net54 _02382_ _02515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06990_ _03198_ _00818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14099_ _01138_ clknet_leaf_145_clk_i memory\[63\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_107_clk_i_I clknet_5_23__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09547__I0 _04631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input7_I data_i[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08660_ _04134_ _01552_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_53_Left_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_89_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07611_ _03209_ memory\[0\]\[27\] _03552_ _03560_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_1_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12059__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08591_ _04097_ _01520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11106__I0 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_72_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07999__I _03751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_124_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_163_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13351__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07542_ memory\[59\]\[27\] _03365_ _03515_ _03523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_92_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07473_ _03485_ _01014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_615 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_9_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_57_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09212_ _04203_ memory\[31\]\[10\] _04441_ _04442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_17_602 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13559__A1 _02902_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_16_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09143_ _04393_ _04405_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08286__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_8_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_44_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11250__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_62_Left_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09719__I _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__A3 _05766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09074_ _04368_ _01732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_47_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_112_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_1047 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08025_ _03790_ _01261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_141_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_40_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07410__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09976_ _04577_ memory\[42\]\[1\] _04861_ _04863_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09538__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12917__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08927_ _04191_ memory\[27\]\[4\] _04286_ _04291_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12298__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_71_Left_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__08210__I0 _03756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08858_ _04254_ _01630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07809_ _03665_ _01170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08789_ _04208_ memory\[25\]\[12\] _04204_ _04209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11425__S _05638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10820_ _05324_ _00442_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_49_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_309_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12470__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10751_ _05070_ memory\[52\]\[31\] _05253_ _05288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13640__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_45_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_109_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13470_ memory\[32\]\[28\] memory\[33\]\[28\] memory\[34\]\[28\] memory\[35\]\[28\]
+ _05670_ _02345_ _02860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_153_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10682_ _05251_ _00377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_36_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_36_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_80_Left_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12421_ _06624_ _00743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_62_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_124_128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11160__S _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10084__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_560 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_35_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15140_ _00099_ clknet_leaf_442_clk_i memory\[43\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12352_ _06555_ _06556_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_69_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11303_ memory\[61\]\[1\] _03128_ _05580_ _05582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15071_ _00030_ clknet_leaf_439_clk_i memory\[41\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12283_ _06467_ _06475_ _06488_ _06489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
Xclkbuf_leaf_284_clk_i clknet_5_14__leaf_clk_i clknet_leaf_284_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_120_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14022_ _01061_ clknet_leaf_247_clk_i memory\[0\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09565__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11234_ _03311_ memory\[60\]\[1\] _05543_ _05545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13595__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12081__S0 _06010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06988__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_140_1050 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_8_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11165_ _05508_ _00603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_8_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_101_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09529__I0 _04619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10116_ _04581_ memory\[44\]\[3\] _04933_ _04937_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_299_clk_i clknet_5_14__leaf_clk_i clknet_leaf_299_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11096_ _03303_ memory\[58\]\[0\] _05471_ _05472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12004__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10047_ _04900_ _00093_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14924_ _01963_ clknet_leaf_48_clk_i memory\[36\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13581__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08909__S _04272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_69_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_89_137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_106_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14855_ _01894_ clknet_leaf_50_clk_i memory\[34\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_222_clk_i clknet_5_26__leaf_clk_i clknet_leaf_222_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_193_4102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13806_ _00845_ clknet_leaf_194_clk_i memory\[16\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_187_356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14786_ _01825_ clknet_leaf_402_clk_i memory\[32\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11998_ _06154_ _06173_ _06190_ _06207_ _06208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__09701__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13737_ _03100_ _00785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_557 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11895__S0 _05742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10949_ _05393_ _00502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_129_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_445 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_237_clk_i clknet_5_26__leaf_clk_i clknet_leaf_237_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_155_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13668_ _05676_ _03050_ _03052_ _03054_ _03055_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_183_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13636__S1 _05726_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12674__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_304 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_827 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15407_ _00366_ clknet_leaf_256_clk_i memory\[51\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12619_ _06467_ _06812_ _06819_ _06820_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__08268__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_33_clk_i_I clknet_5_7__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_735 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_27_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12166__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13599_ memory\[44\]\[30\] memory\[45\]\[30\] _05678_ _02987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11070__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_476 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10075__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15338_ _00297_ clknet_leaf_242_clk_i memory\[4\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_147_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_638 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_42_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_101_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_124_662 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15269_ _00228_ clknet_leaf_404_clk_i memory\[47\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_811 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09393__A1 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09830_ memory\[3\]\[30\] _03217_ _04750_ _04784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10414__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06898__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_165_3558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_258_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09761_ _04637_ memory\[38\]\[30\] _04713_ _04747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06973_ _03185_ _00814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_182_3872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_182_3883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08712_ _03781_ memory\[24\]\[14\] _04157_ _04162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13725__S _03086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09692_ _04710_ _02008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_813 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07723__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08643_ _04125_ _01544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12127__S1 _05922_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08574_ _04088_ _01512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA_clkbuf_leaf_310_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_310 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13244__A3 _02622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07525_ memory\[59\]\[19\] _03348_ _03504_ _03514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13460__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08554__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07456_ _03476_ _01006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_584 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11638__S0 _05778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12076__S _06143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07387_ _03438_ _00975_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_161_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09126_ _04396_ _01756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_165_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_32_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_102_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09057_ _04185_ memory\[2\]\[1\] _04358_ _04360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_323 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09385__S _04524_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08008_ _03165_ _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09759__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_102_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08431__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10324__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09959_ _04853_ _00052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__06993__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12970_ _05677_ _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__08729__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output46_I net46 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11921_ _06085_ _06101_ _06116_ _06131_ _06132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__11663__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09931__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_86_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14640_ _01679_ clknet_leaf_97_clk_i memory\[27\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_47_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11852_ _05788_ _06063_ _05792_ _06064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_68_844 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10803_ _05054_ memory\[53\]\[23\] _05312_ _05316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14571_ _01610_ clknet_leaf_187_clk_i memory\[25\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12443__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11783_ _05950_ _05965_ _05980_ _05995_ _05996_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XPHY_EDGE_ROW_109_Left_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_83_814 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13522_ _02910_ _02911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_10734_ _05279_ _00401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08464__S _04023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_858 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13618__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_24_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13453_ memory\[6\]\[28\] memory\[7\]\[28\] _02322_ _02843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10665_ memory\[51\]\[22\] _03193_ _05240_ _05243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12404_ memory\[30\]\[12\] memory\[31\]\[12\] _06193_ _06608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_35_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13384_ memory\[48\]\[27\] memory\[49\]\[27\] memory\[50\]\[27\] memory\[51\]\[27\]
+ _05725_ _05726_ _02775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_180_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10596_ _05052_ memory\[50\]\[22\] _05203_ _05206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15123_ _00082_ clknet_leaf_11_clk_i memory\[42\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12335_ memory\[30\]\[11\] memory\[31\]\[11\] _06193_ _06540_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07808__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15054_ _00013_ clknet_leaf_20_clk_i memory\[40\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12266_ _05669_ _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XPHY_EDGE_ROW_118_Left_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_82_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_121_687 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_147_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14005_ _01044_ clknet_leaf_160_clk_i memory\[59\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11217_ _05535_ _00628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08422__I0 _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10234__S _04991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput70 net70 data_o[8] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_12197_ _05788_ _06403_ _05792_ _06404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_11148_ _03361_ memory\[58\]\[25\] _05493_ _05499_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11079_ _05462_ _00563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_161_clk_i clknet_5_24__leaf_clk_i clknet_leaf_161_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_160_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_160_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09922__I0 _04591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14907_ _01946_ clknet_leaf_1_clk_i memory\[35\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_37_1035 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11065__S _05446_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_77_129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14838_ _01877_ clknet_leaf_72_clk_i memory\[33\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_127_Left_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_53_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12434__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14769_ _01808_ clknet_leaf_91_clk_i memory\[31\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_176_clk_i clknet_5_28__leaf_clk_i clknet_leaf_176_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_58_365 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07310_ _03397_ _00939_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_128_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10296__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_58_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08290_ _03768_ memory\[18\]\[8\] _03929_ _03938_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07161__I0 _03215_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07241_ _03193_ _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_143_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10048__I0 _04581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07172_ _03307_ _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_119_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_147_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__I1 _03357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_136_Left_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_44_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1197 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11748__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_114_clk_i clknet_5_23__leaf_clk_i clknet_leaf_114_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_111_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_184_3923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_22_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__10220__I0 _04616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09813_ _04775_ _02064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09933__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_696 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_129_clk_i clknet_5_23__leaf_clk_i clknet_leaf_129_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09744_ _04738_ _02032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06956_ _03172_ memory\[14\]\[15\] _03157_ _03173_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_158_1163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07453__S _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13465__A3 _02854_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09675_ _04619_ memory\[37\]\[21\] _04700_ _04702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06887_ net1 _03119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08626_ _04116_ _01536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08557_ _04079_ _01504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12425__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10287__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07508_ _03505_ _01029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12520__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08284__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08488_ _03762_ memory\[21\]\[5\] _04037_ _04043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07439_ memory\[49\]\[11\] _03332_ _03466_ _03468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10450_ _05128_ _00268_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_162_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09109_ _04237_ memory\[2\]\[26\] _04380_ _04387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_60_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10381_ _05041_ memory\[47\]\[17\] _05084_ _05092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12534__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07455__I1 _03348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12120_ _06325_ _06327_ _06328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__07628__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_440 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10054__S _04897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12051_ _05921_ _06259_ _06260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__08404__I0 _03814_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11002_ _05047_ memory\[56\]\[20\] _05421_ _05422_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10211__I0 _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10989__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15810_ _00769_ clknet_leaf_302_clk_i memory\[9\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12489__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15741_ _00700_ clknet_leaf_312_clk_i memory\[62\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_77_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12953_ memory\[46\]\[20\] memory\[47\]\[20\] _06596_ _02351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_93_clk_i clknet_5_20__leaf_clk_i clknet_leaf_93_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_11904_ _05748_ _06110_ _06112_ _06114_ _06115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XTAP_TAPCELL_ROW_29_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15672_ _00631_ clknet_leaf_152_clk_i memory\[5\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12884_ _02209_ _02278_ _02280_ _02282_ _02283_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_73_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_184_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_169_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14623_ _01662_ clknet_leaf_415_clk_i memory\[27\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11835_ memory\[46\]\[4\] memory\[47\]\[4\] _05907_ _06047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12709__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_206_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11613__S _05720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_808 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_28_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10278__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_83_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12967__A2 _02364_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14554_ _01593_ clknet_leaf_3_clk_i memory\[24\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08194__S _03879_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11766_ _05748_ _05974_ _05976_ _05978_ _05979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__07143__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13505_ _05700_ _02889_ _02891_ _02893_ _02894_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__13113__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10717_ _05270_ _00393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_113_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14485_ _01524_ clknet_leaf_105_clk_i memory\[22\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_125_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11697_ _05760_ _05910_ _05911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_153_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_125_245 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_70_327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_82_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13436_ memory\[60\]\[28\] memory\[61\]\[28\] _05702_ _02826_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_733 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_67_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10648_ memory\[51\]\[14\] _03168_ _05229_ _05234_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_183_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_1207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_107_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1327 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_12_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_clk_i clknet_5_7__leaf_clk_i clknet_leaf_31_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_13367_ _02375_ _02758_ _02759_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12444__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10579_ _05035_ memory\[50\]\[14\] _05192_ _05197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07538__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15106_ _00065_ clknet_leaf_442_clk_i memory\[42\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_51_596 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12318_ memory\[36\]\[11\] memory\[37\]\[11\] _06447_ _06523_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12027__S0 _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1040 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13298_ _02494_ _02686_ _02688_ _02690_ _02691_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_114_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15037_ _02076_ clknet_leaf_434_clk_i memory\[40\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12249_ memory\[32\]\[10\] memory\[33\]\[10\] memory\[34\]\[10\] memory\[35\]\[10\]
+ _06314_ _06454_ _06455_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_139_68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09753__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_46_clk_i clknet_5_18__leaf_clk_i clknet_leaf_46_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_177_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08369__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07790_ _03655_ _01161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_147_Right_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_64_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09552__I _03214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_190_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_78 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09460_ _04572_ _01914_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_98 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08411_ _04002_ _01435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09391_ _04247_ memory\[33\]\[31\] _04501_ _04536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_148_337 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_2_2_0_clk_i_I clknet_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_87_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_171_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08342_ _03746_ memory\[1\]\[0\] _03965_ _03966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13080__A1 _06713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07134__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_900 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_75 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_58_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08273_ _03928_ _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10139__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08882__I0 _04214_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_543 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07224_ _03343_ _00907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08832__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_15_755 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_42_541 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07155_ _03206_ memory\[13\]\[26\] _03290_ _03297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12354__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_14_243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07437__I1 _03329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_408_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10441__I0 _05033_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07086_ _03209_ memory\[16\]\[27\] _03251_ _03259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_112_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_974 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07247__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06948__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_2_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_155_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13518__S0 _05784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10602__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07988_ _03765_ _01249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07183__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_114_Right_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09727_ _04729_ _02024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06939_ _03159_ _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__13694__I0 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_9_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12741__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09658_ _04602_ memory\[37\]\[13\] _04689_ _04693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07373__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08609_ _04106_ _01529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_166_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09589_ _04656_ _01959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11433__S _05615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11620_ _05834_ _05835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_93_931 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13071__A1 _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08806__I _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11551_ _03224_ _05767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_53_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09838__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_108_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10502_ _05144_ _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_14270_ _01309_ clknet_leaf_354_clk_i memory\[29\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11482_ _05651_ _05674_ _05697_ _05698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__12257__S0 _06186_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_513 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13221_ memory\[44\]\[24\] memory\[45\]\[24\] _02210_ _02615_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_162_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07428__I1 _03321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_33_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10433_ _05119_ _00260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12264__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_104_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10432__I0 _05024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__S _03415_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13152_ _02546_ _02547_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_131_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10364_ _05024_ memory\[47\]\[9\] _05073_ _05083_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_12103_ _06310_ _06311_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_104_1213 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_20_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13083_ _02478_ _02479_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_130_292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10295_ _03174_ _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09573__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12034_ _05736_ _06242_ _06177_ _06243_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_72_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12885__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__06996__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_137_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12637__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13985_ _01024_ clknet_leaf_324_clk_i memory\[59\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10311__I _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12936_ _06713_ _02329_ _02331_ _02333_ _02334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_15724_ _00683_ clknet_leaf_245_clk_i memory\[61\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_73_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12867_ memory\[8\]\[19\] memory\[9\]\[19\] memory\[10\]\[19\] memory\[11\]\[19\]
+ _06582_ _06721_ _02266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__12439__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15655_ _00614_ clknet_leaf_242_clk_i memory\[5\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11343__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_357_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14606_ _01645_ clknet_leaf_125_clk_i memory\[26\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_68_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11818_ _06028_ _06029_ _05722_ _06030_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_15586_ _00545_ clknet_leaf_319_clk_i memory\[57\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12798_ _06720_ _02197_ _02198_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_185_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_55_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14537_ _01576_ clknet_leaf_174_clk_i memory\[24\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_155_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_155_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11749_ memory\[8\]\[3\] memory\[9\]\[3\] memory\[10\]\[3\] memory\[11\]\[3\] _05893_
+ _05726_ _05962_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_154_852 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_705 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14468_ _01507_ clknet_leaf_363_clk_i memory\[22\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_55_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_116_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_154_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13419_ _02809_ _02810_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_10_1082 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_109_1124 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12174__S _06039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14399_ _01438_ clknet_leaf_353_clk_i memory\[20\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_49_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_51_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_1146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08451__I _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08960_ _04285_ _04308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12902__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07911_ _03719_ _01218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09041__I0 _04237_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08891_ _04271_ _01646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11518__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10422__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07842_ _03147_ memory\[7\]\[7\] _03675_ _03683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08099__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07773_ _03646_ _01153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_179_3811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_179_3822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09512_ _03174_ _04608_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07731__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09443_ _04231_ memory\[34\]\[23\] _04560_ _04564_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12349__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11253__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_611 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09374_ _04527_ _01873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07107__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_192_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_75_964 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08325_ _03956_ _01395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_117_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12800__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08855__I0 _04187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_7_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_10_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09658__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08256_ _03802_ memory\[17\]\[24\] _03915_ _03920_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_81_clk_i_I clknet_5_20__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08562__S _04073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_172_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07207_ _03159_ _03332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_90_989 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_144_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10891__I _05362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08187_ _03883_ _01330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11367__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10414__I0 _05004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07138_ _03181_ memory\[13\]\[18\] _03279_ _03288_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09280__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_37_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_93_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07069_ _03184_ memory\[16\]\[19\] _03240_ _03250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07906__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_54_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10080_ _04917_ _00109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07594__I0 _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12619__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13770_ _00809_ clknet_leaf_201_clk_i memory\[14\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08737__S _04168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10982_ _05411_ _00517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07346__I0 _03129_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12721_ _06844_ _02117_ _02119_ _02121_ _02122_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_139_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11671__B _05708_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_955 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_97_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15440_ _00399_ clknet_leaf_261_clk_i memory\[52\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12652_ memory\[0\]\[16\] memory\[1\]\[16\] memory\[2\]\[16\] memory\[3\]\[16\] _06709_
+ _06779_ _06852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09099__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13044__A1 _02375_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12478__S0 _06342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_154_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11603_ _05651_ _05810_ _05817_ _05818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_33_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_182_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15371_ _00330_ clknet_leaf_240_clk_i memory\[50\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12583_ _06783_ _06784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_26_828 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_81_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14322_ _01361_ clknet_leaf_103_clk_i memory\[17\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_92_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11534_ memory\[44\]\[0\] memory\[45\]\[0\] _05749_ _05750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08472__S _04000_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_14253_ _01292_ clknet_leaf_199_clk_i memory\[15\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11465_ _03118_ _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10507__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_179 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07088__S _03251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13204_ _06851_ _02597_ _02598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_151_888 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10416_ _05008_ memory\[48\]\[1\] _05109_ _05111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14184_ _01223_ clknet_leaf_206_clk_i memory\[19\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09271__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11396_ _03336_ memory\[62\]\[13\] _05627_ _05631_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_74_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10956__I1 _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_81_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_111_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13135_ _02302_ _02522_ _02529_ _02530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XTAP_TAPCELL_ROW_111_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12722__S _06714_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10347_ _05074_ _00219_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_108_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07816__S _03661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13066_ memory\[4\]\[22\] memory\[5\]\[22\] _06845_ _02462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10278_ _05026_ memory\[46\]\[10\] _05027_ _05028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11338__S _05591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12017_ _06225_ _06226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_139_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10242__S _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11530__A1 _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_174_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13553__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11137__I _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10041__I _04896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13968_ _01007_ clknet_leaf_161_clk_i memory\[49\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_15707_ _00666_ clknet_leaf_389_clk_i memory\[60\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_157_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12919_ _06831_ _02311_ _02314_ _02316_ _02317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_186_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13899_ _00938_ clknet_leaf_209_clk_i memory\[11\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_0_36 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_100_Left_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_186_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_158_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13035__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15638_ _00597_ clknet_leaf_160_clk_i memory\[58\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_174_3730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_8_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_173_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_84_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_189_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_103_clk_i_I clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15569_ _00528_ clknet_leaf_169_clk_i memory\[56\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_08110_ _03793_ memory\[15\]\[20\] _03841_ _03842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_170_3649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09090_ _04218_ memory\[2\]\[17\] _04369_ _04377_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_154_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_4_711 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08041_ _03801_ _01266_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_25_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_395 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09992_ _04593_ memory\[42\]\[9\] _04861_ _04871_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_52 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09014__I0 _04210_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08943_ _04299_ _01670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11756__B _05739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_983 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_85 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11248__S _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10152__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08874_ _04206_ memory\[26\]\[11\] _04261_ _04263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_32_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07576__I0 _03156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_28_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09941__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07825_ _03673_ _01178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_93_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07756_ _03221_ memory\[63\]\[31\] _03602_ _03637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13274__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09740__I _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07687_ _03600_ _01113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_454 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10883__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09426_ _04214_ memory\[34\]\[15\] _04549_ _04555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_164_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09357_ _04518_ _01865_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_3__f_clk_i clknet_2_0_0_clk_i clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08308_ _03947_ _01387_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08292__S _03929_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09288_ _04212_ memory\[32\]\[14\] _04477_ _04482_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_95_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_133_833 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_95_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08239_ _03785_ memory\[17\]\[16\] _03904_ _03911_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_593 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_132_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_65_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10327__S _05048_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11510__I _05693_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_820 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_132_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11250_ _03327_ memory\[60\]\[9\] _05543_ _05553_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09253__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_91_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_120_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10938__I1 _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_305_clk_i_I clknet_5_11__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10201_ _04598_ memory\[45\]\[11\] _04980_ _04982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12542__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11181_ _05516_ _00611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_101_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07636__S _03567_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10132_ _04945_ _00133_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13188__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09005__I0 _04201_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_100_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_1276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11158__S _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14940_ _01979_ clknet_leaf_435_clk_i memory\[37\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10063_ _04595_ memory\[43\]\[10\] _04908_ _04909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07567__I0 _03144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11512__A1 _05724_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11363__I1 _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14871_ _01910_ clknet_leaf_73_clk_i memory\[34\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10997__S _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13373__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_1041 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13822_ _00861_ clknet_leaf_373_clk_i memory\[13\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_173_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13265__A1 _06848_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_134_1014 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07371__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13753_ _03108_ _00793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10796__I _05289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10965_ _05402_ _00509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_1069 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12704_ memory\[56\]\[17\] memory\[57\]\[17\] memory\[58\]\[17\] memory\[59\]\[17\]
+ _06827_ _06280_ _02105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_57_227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_67_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_67_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13684_ _03224_ _03063_ _03070_ _03071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_104_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10896_ memory\[55\]\[2\] _03131_ _05363_ _05366_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_191_4052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_155_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_122_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15423_ _00382_ clknet_leaf_331_clk_i memory\[52\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12635_ _05681_ _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_54_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12717__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11621__S _05737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_794 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09298__S _04477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_53_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15354_ _00313_ clknet_leaf_392_clk_i memory\[4\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_142_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12566_ memory\[52\]\[15\] memory\[53\]\[15\] _06143_ _06767_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_170_438 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14305_ _01344_ clknet_leaf_344_clk_i memory\[17\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11517_ _05655_ _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_15285_ _00244_ clknet_leaf_385_clk_i memory\[47\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_135_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_628 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12497_ _05691_ _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_0_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14236_ _01275_ clknet_leaf_278_clk_i memory\[15\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11448_ _03112_ _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_141_1007 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_33_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__10929__I1 _03180_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11051__I0 _05029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14167_ _01206_ clknet_leaf_140_clk_i memory\[7\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09795__I1 _03165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12452__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11379_ _03319_ memory\[62\]\[5\] _05616_ _05622_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11751__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07546__S _03515_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13118_ _02461_ _02477_ _02493_ _02513_ _02514_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_0_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14098_ _01137_ clknet_leaf_133_clk_i memory\[63\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13049_ _02445_ _00752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09761__S _04713_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07610_ _03559_ _01077_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_1_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08590_ _03796_ memory\[22\]\[21\] _04095_ _04097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08377__S _03976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_124_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_178_549 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07541_ _03522_ _01045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13351__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_763 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10865__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13008__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07472_ memory\[49\]\[27\] _03365_ _03477_ _03485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09211_ _04429_ _04441_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_147_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_435 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13559__A2 _02917_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_254_clk_i_I clknet_5_24__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_45_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_5_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_405_clk_i clknet_5_3__leaf_clk_i clknet_leaf_405_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_934 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_17_636 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09142_ _04404_ _01764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_72_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_45_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09001__S _04322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09073_ _04201_ memory\[2\]\[9\] _04358_ _04368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11290__I0 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11585__A4 _05800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10147__S _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08024_ _03789_ memory\[12\]\[18\] _03773_ _03790_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09235__I0 _04227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_40 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13458__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11042__I0 _05020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__I1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_187_3965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07797__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09975_ _04862_ _00059_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07410__A2 net6 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08926_ _04290_ _01662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12917__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13495__A1 _02358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11345__I1 _03190_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_157_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08857_ _04189_ memory\[26\]\[3\] _04250_ _04254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13193__S _02312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07808_ _03197_ memory\[6\]\[23\] _03661_ _03665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_100_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10610__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08788_ _03162_ _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_79_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07739_ _03628_ _01137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_49_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10856__I0 _05039_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10750_ _05287_ _00409_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_177_582 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07721__I0 _03169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09409_ _04197_ memory\[34\]\[7\] _04538_ _04546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_295 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10681_ memory\[51\]\[30\] _03217_ _05217_ _05251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11441__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10608__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12420_ _06623_ net43 _06491_ _06624_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_152_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_36_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_62_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12351_ memory\[60\]\[12\] memory\[61\]\[12\] _06273_ _06555_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_129_1149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_11302_ _05581_ _00667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09846__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_121_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15070_ _00029_ clknet_leaf_440_clk_i memory\[41\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09226__I0 _04218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12282_ _06476_ _06479_ _06483_ _06487_ _06488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_15_190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14021_ _01060_ clknet_leaf_338_clk_i memory\[0\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_31_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11233_ _05544_ _00635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_120_335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12272__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11733__A1 _05682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12081__S1 _06150_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_30_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11164_ _03303_ memory\[5\]\[0\] _05507_ _05508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_8_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_105_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10115_ _04936_ _00125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12071__I _05667_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13486__A1 _02501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11095_ _05470_ _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_175_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11336__I1 _03177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09581__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_145_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10046_ _04579_ memory\[43\]\[2\] _04897_ _04900_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14923_ _01962_ clknet_leaf_47_clk_i memory\[36\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13581__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_69_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_69_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14854_ _01893_ clknet_leaf_52_clk_i memory\[34\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_188_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07960__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_193_4114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13805_ _00844_ clknet_leaf_206_clk_i memory\[16\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11997_ _05767_ _06199_ _06206_ _06207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_14785_ _01824_ clknet_leaf_419_clk_i memory\[32\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_97_160 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13736_ _03355_ memory\[9\]\[22\] _03097_ _03100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10948_ memory\[55\]\[27\] _03208_ _05385_ _05393_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_48 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08925__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11895__S1 _05743_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12955__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13667_ _05690_ _03053_ _03054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10879_ _05062_ memory\[54\]\[27\] _05348_ _05356_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_186_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11351__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_720 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_27_945 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_1175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15406_ _00365_ clknet_leaf_259_clk_i memory\[51\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12618_ _06476_ _06814_ _06816_ _06818_ _06819_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08724__I _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_26_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13598_ _05654_ _02981_ _02983_ _02985_ _02986_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_0_109_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12549_ _05701_ _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_136_490 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15337_ _00296_ clknet_leaf_242_clk_i memory\[4\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_391_clk_i clknet_5_3__leaf_clk_i clknet_leaf_391_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_15268_ _00227_ clknet_leaf_405_clk_i memory\[47\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_302 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11024__I0 _05070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14219_ _01258_ clknet_leaf_198_clk_i memory\[12\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09768__I1 _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15199_ _00158_ clknet_leaf_438_clk_i memory\[45\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_10_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09555__I _03217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07276__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09393__A2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13077__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_165_3559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09760_ _04746_ _02040_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06972_ _03184_ memory\[14\]\[19\] _03157_ _03185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13021__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_126_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09491__S _04575_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08711_ _04161_ _01576_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09691_ _04635_ memory\[37\]\[29\] _04700_ _04710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_119_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08642_ memory\[23\]\[13\] _03336_ _04121_ _04125_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10430__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_90_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08573_ _03779_ memory\[22\]\[13\] _04084_ _04088_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07524_ _03513_ _01037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08835__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_344_clk_i clknet_5_8__leaf_clk_i clknet_leaf_344_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_14_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_5_21__f_clk_i clknet_2_2_0_clk_i clknet_5_21__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_130_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_18_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07455_ memory\[49\]\[19\] _03348_ _03466_ _03476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_14_1058 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_162_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11261__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_574 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07386_ _03187_ memory\[8\]\[20\] _03437_ _03438_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13401__A1 _05768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_416 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_106_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11638__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09125_ _04185_ memory\[30\]\[1\] _04394_ _04396_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_44_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11263__I0 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_359_clk_i clknet_5_2__leaf_clk_i clknet_leaf_359_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_33_937 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_40_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11963__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_72_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_161_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09666__S _04689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09056_ _04359_ _01723_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_124_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_130_633 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08007_ _03778_ _01255_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_163_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12092__S _06025_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11715__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07186__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_688 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13180__A3 _02574_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12105__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_5_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09958_ _04627_ memory\[41\]\[25\] _04847_ _04853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07914__S _03711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_95_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08909_ _04241_ memory\[26\]\[28\] _04272_ _04281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09889_ _04816_ _00019_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11920_ _05767_ _06123_ _06130_ _06131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_86_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08809__I _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07942__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11851_ memory\[22\]\[4\] memory\[23\]\[4\] _06062_ _06063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_169_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10829__I0 _05012_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_1250 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10802_ _05315_ _00433_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14570_ _01609_ clknet_leaf_187_clk_i memory\[25\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11782_ _05767_ _05987_ _05994_ _05995_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08745__S _04145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09695__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_390 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13521_ memory\[12\]\[29\] memory\[13\]\[29\] _05769_ _02910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_83_826 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10733_ _05052_ memory\[52\]\[22\] _05276_ _05279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_71_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13452_ _02841_ _02842_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__09447__I0 _04235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10664_ _05242_ _00368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12826__S0 _06472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_82_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12403_ _05659_ _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_106_630 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13383_ _05719_ _02773_ _02178_ _02774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_10595_ _05205_ _00336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_296 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11954__A1 _06162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12334_ _06538_ _06539_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_15122_ _00081_ clknet_leaf_13_clk_i memory\[42\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08480__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_50_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07622__A2 net72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11006__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15053_ _00012_ clknet_leaf_24_clk_i memory\[40\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12265_ _05918_ _06470_ _06195_ _06471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__06999__I net25 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_981 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10515__S _05156_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13251__S0 _06827_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_128_Right_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11706__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14004_ _01043_ clknet_leaf_166_clk_i memory\[59\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11216_ _03361_ memory\[5\]\[25\] _05529_ _05535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_202_clk_i_I clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12196_ memory\[22\]\[9\] memory\[23\]\[9\] _06062_ _06403_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput60 net60 data_o[28] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
Xoutput71 net71 data_o[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_120_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11147_ _05498_ _00595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10314__I _03193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12730__S _06447_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_1317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11309__I1 _03137_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07824__S _03638_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1091 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11078_ _05056_ memory\[57\]\[24\] _05457_ _05462_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08186__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10250__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14906_ _01945_ clknet_leaf_5_clk_i memory\[35\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_10029_ _04890_ _00085_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_160_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07933__I0 _03181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07623__I _03566_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_192_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14837_ _01876_ clknet_leaf_74_clk_i memory\[33\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_121_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_114_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14768_ _01807_ clknet_leaf_90_clk_i memory\[31\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13631__A1 _05700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_85_130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12685__B _02086_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_517 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13719_ _03338_ memory\[9\]\[14\] _03086_ _03091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_18_219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_232 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14699_ _01738_ clknet_leaf_176_clk_i memory\[2\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07240_ _03354_ _00912_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_184_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_6_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07171_ _03305_ _03306_ _03307_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__12905__S _02164_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_119_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08110__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_42_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_419 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08390__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_136_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__06903__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08661__I1 _03355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_124_482 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_78_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_169_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_83_1078 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13736__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12370__A1 _06159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09812_ memory\[3\]\[21\] _03190_ _04773_ _04775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07734__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_06955_ _03171_ _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_09743_ _04619_ memory\[38\]\[21\] _04736_ _04738_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08177__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12122__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10160__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09674_ _04701_ _01999_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06886_ _03116_ _03117_ _03118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_94_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08625_ memory\[23\]\[5\] _03319_ _04110_ _04116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_404_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_283_clk_i clknet_5_14__leaf_clk_i clknet_leaf_283_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_167_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08556_ _03762_ memory\[22\]\[5\] _04073_ _04079_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13622__A1 _02964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09677__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12425__A2 _06627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_92_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07507_ memory\[59\]\[10\] _03329_ _03504_ _03505_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08487_ _04042_ _01471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12087__S _05706_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_42_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_21_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07438_ _03467_ _00997_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_147_585 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_80_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_736 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_151_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_21_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_64_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_298_clk_i clknet_5_14__leaf_clk_i clknet_leaf_298_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_162_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11236__I0 _03313_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07369_ _03163_ memory\[8\]\[12\] _03426_ _03429_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08101__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09108_ _04386_ _01748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10380_ _05091_ _00235_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08652__I1 _03346_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_791 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_221_clk_i clknet_5_27__leaf_clk_i clknet_leaf_221_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_09039_ _04235_ memory\[28\]\[25\] _04344_ _04350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_27_1238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12050_ memory\[24\]\[7\] memory\[25\]\[7\] memory\[26\]\[7\] memory\[27\]\[7\] _05778_
+ _05922_ _06259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_57_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11001_ _05398_ _05421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__12550__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_236_clk_i clknet_5_26__leaf_clk_i clknet_leaf_236_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_142_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11547__S0 _05761_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11166__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15740_ _00699_ clknet_leaf_311_clk_i memory\[62\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_76_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12952_ _02349_ _02350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_176_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_137_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_88_929 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11903_ _05760_ _06113_ _06114_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_59_108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15671_ _00630_ clknet_leaf_151_clk_i memory\[5\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_29_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_38_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_29_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_1247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12883_ _02216_ _02281_ _02282_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_14622_ _01661_ clknet_leaf_415_clk_i memory\[27\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11834_ _06045_ _06046_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__12416__A2 _06619_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_56_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13613__A1 _02494_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09668__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14553_ _01592_ clknet_leaf_78_clk_i memory\[24\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11765_ _05760_ _05977_ _05978_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_138_563 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_55_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13504_ _05710_ _02892_ _02893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_10716_ _05035_ memory\[52\]\[14\] _05265_ _05270_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14484_ _01523_ clknet_leaf_105_clk_i memory\[22\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11696_ memory\[40\]\[2\] memory\[41\]\[2\] memory\[42\]\[2\] memory\[43\]\[2\] _05761_
+ _05762_ _05910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_187_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_70_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10647_ _05233_ _00360_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13435_ _02825_ _00758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_64_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1275 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11927__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13366_ memory\[16\]\[26\] memory\[17\]\[26\] memory\[18\]\[26\] memory\[19\]\[26\]
+ _02233_ _02376_ _02758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_144_1219 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_10578_ _05196_ _00328_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09840__I0 _04577_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15105_ _00064_ clknet_leaf_439_clk_i memory\[42\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_5_29__f_clk_i_I clknet_2_3_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12317_ _06428_ _06514_ _06521_ _06522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_13297_ _02501_ _02689_ _02690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_23_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12027__S1 _06032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_107_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_114_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15036_ _02075_ clknet_leaf_435_clk_i memory\[40\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12248_ _03747_ _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_139_47 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_353_clk_i_I clknet_5_2__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12179_ memory\[44\]\[9\] memory\[45\]\[9\] _06319_ _06386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08159__I0 _03772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11076__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_155_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_79_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_155_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07906__I0 _03141_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_64_77 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08410_ _03746_ memory\[20\]\[0\] _04001_ _04002_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_8_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_118_1181 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09390_ _04535_ _01881_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13604__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_74_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08341_ _03964_ _03965_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_177_3783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_15_1142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_54_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_606 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_168 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_50 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_157_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_149_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08272_ _03225_ net72 _03928_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_07223_ memory\[39\]\[16\] _03342_ _03330_ _03343_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11218__I0 _03363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10219__I _04968_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11918__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_588 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07729__S _03614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07154_ _03296_ _00884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_255 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07085_ _03258_ _00853_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_30_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_113_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13135__A3 _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12343__A1 _06480_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08398__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13466__S _02338_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1203 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07464__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input38_I data_i[9] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13518__S1 _03226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_35_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07987_ _03764_ memory\[12\]\[6\] _03752_ _03765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09726_ _04602_ memory\[38\]\[13\] _04725_ _04729_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06938_ net9 _03159_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__09898__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09657_ _04692_ _01991_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_145_90 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_26_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11714__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_625 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_136_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08608_ _03814_ memory\[22\]\[30\] _04072_ _04106_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08295__S _03940_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09588_ _04600_ memory\[36\]\[12\] _04653_ _04656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_496 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08539_ _04069_ _01496_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08322__I0 _03800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_617 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_38_859 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11550_ _05731_ _05746_ _05765_ _05766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_0_64_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_93_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10501_ _05155_ _00292_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11481_ _05676_ _05680_ _05688_ _05696_ _05697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_190_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11909__A1 _05918_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12257__S1 _06326_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_98_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13220_ _02337_ _02609_ _02611_ _02613_ _02614_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_107_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_160_clk_i clknet_5_25__leaf_clk_i clknet_leaf_160_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_10432_ _05024_ memory\[48\]\[9\] _05109_ _05119_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08822__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08625__I1 _03319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_59_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13151_ memory\[36\]\[23\] memory\[37\]\[23\] _02338_ _02546_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_33_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10363_ _05082_ _00227_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10065__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12102_ memory\[36\]\[8\] memory\[37\]\[8\] _05733_ _06310_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_20_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09854__S _04789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_76_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13082_ memory\[36\]\[22\] memory\[37\]\[22\] _02338_ _02478_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10294_ _05038_ _00202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_175_clk_i clknet_5_28__leaf_clk_i clknet_leaf_175_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12033_ memory\[38\]\[7\] memory\[39\]\[7\] _06039_ _06242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10196__I0 _04593_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_155_Left_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_72_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07061__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_72_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_18_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13984_ _01023_ clknet_leaf_323_clk_i memory\[59\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07173__I _03308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_77_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15723_ _00682_ clknet_leaf_245_clk_i memory\[61\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12935_ _06720_ _02332_ _02333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_0_88_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15654_ _00613_ clknet_leaf_244_clk_i memory\[5\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_115_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12866_ _06717_ _02264_ _02195_ _02265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
Xclkbuf_leaf_113_clk_i clknet_5_23__leaf_clk_i clknet_leaf_113_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_14605_ _01644_ clknet_leaf_124_clk_i memory\[26\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12519__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13124__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_837 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11817_ memory\[14\]\[4\] memory\[15\]\[4\] _05720_ _06029_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_157_157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15585_ _00544_ clknet_5_10__leaf_clk_i memory\[57\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_185_477 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08313__I0 _03791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12797_ memory\[8\]\[18\] memory\[9\]\[18\] memory\[10\]\[18\] memory\[11\]\[18\]
+ _06582_ _06721_ _02197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_164_Left_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_28_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11999__I1 net68 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14536_ _01575_ clknet_leaf_183_clk_i memory\[24\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08933__S _04286_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10120__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11748_ _05719_ _05960_ _05722_ _05961_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_155_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_382 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_12_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10671__I1 _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14467_ _01506_ clknet_leaf_350_clk_i memory\[22\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11679_ _05691_ _05893_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_TAPCELL_ROW_116_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_128_clk_i clknet_5_23__leaf_clk_i clknet_leaf_128_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_172_3691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_181_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13418_ memory\[28\]\[27\] memory\[29\]\[27\] _02495_ _02809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_144_1005 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14398_ _01437_ clknet_leaf_352_clk_i memory\[20\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_180_Right_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_133_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12573__A1 _06411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_249 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13349_ memory\[46\]\[26\] memory\[47\]\[26\] _02487_ _02741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_59_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13117__A3 _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_173_Left_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__13286__S _02487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15019_ _02058_ clknet_leaf_170_clk_i memory\[3\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_07910_ _03147_ memory\[19\]\[7\] _03711_ _03719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_08890_ _04222_ memory\[26\]\[19\] _04261_ _04271_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10703__S _05254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12876__A2 _02274_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07284__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07841_ _03682_ _01185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_75_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10502__I _05144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08179__I _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07772_ _03144_ memory\[6\]\[6\] _03639_ _03646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_79_704 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09511_ _04607_ _01930_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_179_3823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_116_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_189_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08552__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11534__S _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_78_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09442_ _04563_ _01905_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_188_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_182_Left_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09373_ _04229_ memory\[33\]\[22\] _04524_ _04527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09257__A1 net73 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_634 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_191_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08324_ _03802_ memory\[18\]\[24\] _03951_ _03956_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_117_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_46_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09939__S _04836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_19_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_998 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08255_ _03919_ _01362_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_24_clk_i_I clknet_5_4__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_89_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07206_ _03331_ _00901_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_6_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08186_ _03800_ memory\[29\]\[23\] _03879_ _03883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_558 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11367__A2 _03490_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12564__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07137_ _03287_ _00876_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_92_clk_i clknet_5_21__leaf_clk_i clknet_leaf_92_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_28_1355 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_191_Left_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_37_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07068_ _03249_ _00845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12316__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10178__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_249_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13209__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11508__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_96_1055 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_57_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09709_ _04585_ memory\[38\]\[5\] _04714_ _04720_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_173_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_69_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10981_ _05026_ memory\[56\]\[10\] _05410_ _05411_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_30_clk_i clknet_5_6__leaf_clk_i clknet_leaf_30_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_179_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12720_ _06851_ _02120_ _02121_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_35_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_70_1217 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10350__I0 _05010_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_301_clk_i_I clknet_5_14__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_38_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_78_781 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12651_ _03117_ _06851_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_182_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12478__S1 _06485_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_137_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11602_ _05676_ _05812_ _05814_ _05816_ _05817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_12582_ memory\[12\]\[15\] memory\[13\]\[15\] _06714_ _06783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_38_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10102__I0 _04635_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15370_ _00329_ clknet_leaf_238_clk_i memory\[50\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_108_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_45_clk_i clknet_5_18__leaf_clk_i clknet_leaf_45_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_68_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14321_ _01360_ clknet_leaf_117_clk_i memory\[17\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_170_609 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12275__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11533_ _05677_ _05749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_108_555 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_135_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_108_577 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07369__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14252_ _01291_ clknet_leaf_199_clk_i memory\[15\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11464_ _05679_ _05680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_34_873 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12555__A1 _06467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_150_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13203_ memory\[0\]\[24\] memory\[1\]\[24\] memory\[2\]\[24\] memory\[3\]\[24\] _05784_
+ _06779_ _02597_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_10415_ _05110_ _00251_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_21_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14183_ _01222_ clknet_leaf_202_clk_i memory\[19\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11395_ _05630_ _00711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_81_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_406 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_21_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09584__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_111_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10346_ _05004_ memory\[47\]\[0\] _05073_ _05074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_271 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13134_ _06831_ _02524_ _02526_ _02528_ _02529_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_103_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11619__S _05733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13065_ _02302_ _02453_ _02460_ _02461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_40_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_1021 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10277_ _05005_ _05027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07034__I0 _03132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12016_ memory\[4\]\[7\] memory\[5\]\[7\] _06156_ _06225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_40_1076 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11530__A2 _05735_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_79_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_26 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_136_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07832__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_501 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12958__B _02353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_109_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_191_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13967_ _01006_ clknet_leaf_242_clk_i memory\[49\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08534__I0 _03808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15706_ _00665_ clknet_leaf_379_clk_i memory\[60\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_567 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12918_ _06838_ _02315_ _02316_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_9_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13898_ _00937_ clknet_leaf_213_clk_i memory\[11\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_157_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_29_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15637_ _00596_ clknet_leaf_160_clk_i memory\[58\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_174_3720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_158_466 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10892__I1 _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12849_ _02247_ _02248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_111_1004 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1173 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13666__S0 _05692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_186_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_5_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_442 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09759__S _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08663__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15568_ _00527_ clknet_leaf_176_clk_i memory\[56\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_28_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_16_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_84_795 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14519_ _01558_ clknet_leaf_105_clk_i memory\[23\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_497 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10644__I1 _03162_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_170_3639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_142_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15499_ _00458_ clknet_leaf_240_clk_i memory\[54\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_43_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_86_1246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08040_ _03800_ memory\[12\]\[23\] _03794_ _03801_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_198_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09558__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12546__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_821 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__06911__S _03126_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_12_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09991_ _04870_ _00067_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_951 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08942_ _04206_ memory\[27\]\[11\] _04297_ _04299_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_250_clk_i_I clknet_5_25__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08873_ _04262_ _01637_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_32_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13744__S _03097_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08773__I0 _04197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07824_ _03221_ memory\[6\]\[31\] _03638_ _03673_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08838__S _04225_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07742__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_07755_ _03636_ _01145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07328__I1 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07686_ _03218_ memory\[10\]\[30\] _03566_ _03600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09425_ _04554_ _01897_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_17_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_109_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08573__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09356_ _04212_ memory\[33\]\[14\] _04513_ _04518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_136_149 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08307_ _03785_ memory\[18\]\[16\] _03940_ _03947_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10635__I1 _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12095__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09287_ _04481_ _01832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_133_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10608__S _05203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_133_823 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07189__S _03309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07500__I1 _03323_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08238_ _03910_ _01354_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_95_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_95_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_62_478 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12537__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_43_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08169_ _03783_ memory\[29\]\[15\] _03868_ _03874_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_31_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_43_692 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10200_ _04981_ _00165_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07917__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11180_ _03325_ memory\[5\]\[8\] _05507_ _05516_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_24_1038 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10131_ _04595_ memory\[44\]\[10\] _04944_ _04945_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output69_I net69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10062_ _04896_ _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__08764__I0 _04191_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11512__A2 _05727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14870_ _01909_ clknet_leaf_72_clk_i memory\[34\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10571__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13821_ _00860_ clknet_leaf_270_clk_i memory\[13\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11174__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_707 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13752_ _03371_ memory\[9\]\[30\] _03074_ _03108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_168_731 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10964_ _05010_ memory\[56\]\[2\] _05399_ _05402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_70_1003 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_887 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_156_904 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12703_ _06276_ _02103_ _06690_ _02104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_70_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13683_ _05748_ _03065_ _03067_ _03069_ _03070_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_TAPCELL_ROW_67_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_712 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_403 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10895_ _05365_ _00476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_104_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_167_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_127_105 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_1335 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15422_ _00381_ clknet_leaf_346_clk_i memory\[52\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09579__S _04642_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_156_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12634_ _06833_ _06834_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_182_244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_152_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_152_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_93_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15353_ _00312_ clknet_leaf_152_clk_i memory\[4\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_81_743 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12565_ _06272_ _06761_ _06763_ _06765_ _06766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__11701__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14304_ _01343_ clknet_leaf_349_clk_i memory\[17\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11516_ _05653_ _05732_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_80_253 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15284_ _00243_ clknet_leaf_39_clk_i memory\[47\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12496_ _06146_ _06697_ _06287_ _06698_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12528__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14235_ _01274_ clknet_leaf_394_clk_i memory\[12\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_80_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10317__I _03196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_139 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11447_ memory\[62\]\[0\] memory\[63\]\[0\] _05662_ _05663_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_85_1290 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_111_528 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14166_ _01205_ clknet_leaf_141_clk_i memory\[7\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11378_ _05621_ _00703_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11349__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13117_ _02358_ _02505_ _02512_ _02513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_10329_ _03208_ _05062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10253__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14097_ _01136_ clknet_leaf_133_clk_i memory\[63\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12387__S0 _06314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_167_3590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13048_ _02444_ net53 _02382_ _02445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_56_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08755__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13564__S _02448_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10562__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11592__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08507__I0 _03781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14999_ _02038_ clknet_leaf_18_clk_i memory\[38\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11084__S _05457_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_178_539 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07540_ memory\[59\]\[26\] _03363_ _03515_ _03522_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_353 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_1261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_152_1137 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_1268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07471_ _03484_ _01013_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_159_797 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1043 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09210_ _04440_ _01796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_118_116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13559__A3 _02932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_146_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09141_ _04201_ memory\[30\]\[9\] _04394_ _04404_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10428__S _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_979 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_694 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09072_ _04367_ _01731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_60_938 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_653 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08023_ _03180_ _03789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_47_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_25_1325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_364 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_40_673 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11259__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09974_ _04573_ memory\[42\]\[0\] _04861_ _04862_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09952__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08925_ _04189_ memory\[27\]\[3\] _04286_ _04290_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_23_1093 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08856_ _04253_ _01629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_157_1048 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_99_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input20_I data_i[21] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07472__S _03477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_80 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07807_ _03664_ _01169_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_19_1107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08787_ _04207_ _01606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_88_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_135_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07738_ _03194_ memory\[63\]\[22\] _03625_ _03628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10305__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_39_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_49_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09171__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_509 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07669_ _03591_ _01104_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_926 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_274 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09399__S _04538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09408_ _04545_ _01889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10680_ _05250_ _00376_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09339_ _04195_ memory\[33\]\[6\] _04502_ _04509_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_109_Right_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__11521__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_62_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_192_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_180_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_129_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_62_231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_164_1008 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_1128 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12350_ _06554_ _00742_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_11301_ memory\[61\]\[0\] _03110_ _05580_ _05581_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13649__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12281_ _06484_ _06486_ _06487_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_160_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_50_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_50_459 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07647__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11232_ _03303_ memory\[60\]\[0\] _05543_ _05544_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14020_ _01059_ clknet_leaf_369_clk_i memory\[0\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09926__I _04824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11163_ _05506_ _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA__10073__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10792__I0 _05043_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10114_ _04579_ memory\[44\]\[2\] _04933_ _04936_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_101_583 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_8_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11094_ _03490_ _03565_ _05470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_179_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__08737__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_175_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_146_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10045_ _04899_ _00092_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11497__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14922_ _01961_ clknet_leaf_35_clk_i memory\[36\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10801__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08478__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10544__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_69_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14853_ _01892_ clknet_leaf_400_clk_i memory\[34\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_106_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_193_4104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13804_ _00843_ clknet_leaf_193_clk_i memory\[16\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_193_4115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14784_ _01823_ clknet_leaf_418_clk_i memory\[32\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11996_ _05783_ _06201_ _06203_ _06205_ _06206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_187_358 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09162__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12997__A1 _06835_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13735_ _03099_ _00784_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10947_ _05392_ _00501_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_58_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_151_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13666_ memory\[40\]\[31\] memory\[41\]\[31\] memory\[42\]\[31\] memory\[43\]\[31\]
+ _05692_ _05694_ _03053_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_156_756 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10878_ _05355_ _00469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_2_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_15405_ _00364_ clknet_leaf_257_clk_i memory\[51\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_183_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12617_ _06484_ _06817_ _06818_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_27_957 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_586 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13597_ _05668_ _02984_ _02985_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_143_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15336_ _00295_ clknet_leaf_238_clk_i memory\[4\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12548_ _06749_ _06750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_170_236 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_170_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_54_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_1216 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_973 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_124_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_112_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15267_ _00226_ clknet_leaf_411_clk_i memory\[47\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_112_815 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12479_ _06484_ _06681_ _06682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_169_3630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07557__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14218_ _01257_ clknet_leaf_202_clk_i memory\[12\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15198_ _00157_ clknet_leaf_438_clk_i memory\[45\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_111_347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_846 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_10_857 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14149_ _01188_ clknet_leaf_294_clk_i memory\[7\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_191_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_165_3549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09772__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06971_ _03183_ _03184_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__13021__S1 _02345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13294__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08710_ _03779_ memory\[24\]\[13\] _04157_ _04161_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13721__I0 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_193_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_TAPCELL_ROW_182_3885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08388__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09690_ _04709_ _02007_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_174_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07292__S _03379_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07400__I0 _03209_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08641_ _04124_ _01543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12780__S0 _06699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_55_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_1032 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08572_ _04087_ _01511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_107_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07523_ memory\[59\]\[18\] _03346_ _03504_ _03513_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_88_194 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_414 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_348_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_159_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07454_ _03475_ _01005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_135_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09012__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_18_935 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13042__B _02373_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_9_678 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_44_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07385_ _03414_ _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_147_789 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_128_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10158__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_726 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_146_277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1287 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08408__A2 _03750_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_161_214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_96_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_134_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09124_ _04395_ _01755_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08851__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12881__B _06461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09055_ _04181_ memory\[2\]\[0\] _04358_ _04359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_128_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_400_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_163_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13165__A1 _02336_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08006_ _03777_ memory\[12\]\[12\] _03773_ _03778_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_41_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_124_1025 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08967__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_60_1046 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_21_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_25_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_5_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09957_ _04852_ _00051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_5_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08908_ _04280_ _01654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10621__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10526__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09888_ _04625_ memory\[40\]\[24\] _04811_ _04816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09481__I _03143_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08839_ _04242_ _01623_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13217__B _06866_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11516__I _05653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_802 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11850_ _05701_ _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_135_1132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_170_1023 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_140_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09144__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_79_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10801_ _05052_ memory\[53\]\[22\] _05312_ _05315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_95_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11781_ _05783_ _05989_ _05991_ _05993_ _05994_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_64_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13731__I _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_101_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_339 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_138_734 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13520_ _05747_ _02904_ _02906_ _02908_ _02909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_101_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10732_ _05278_ _00400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08825__I _03199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_531 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13451_ memory\[4\]\[28\] memory\[5\]\[28\] _05789_ _02841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10663_ memory\[51\]\[21\] _03190_ _05240_ _05242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12826__S1 _06611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12402_ _06605_ _06606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_137_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_439 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08761__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13382_ memory\[54\]\[27\] memory\[55\]\[27\] _02312_ _02773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10594_ _05050_ memory\[50\]\[21\] _05203_ _05205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_72_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15121_ _00080_ clknet_leaf_7_clk_i memory\[42\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_90_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12333_ memory\[28\]\[11\] memory\[29\]\[11\] _05915_ _06538_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_133_450 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_19__f_clk_i_I clknet_2_2_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_675 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07377__S _03426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15052_ _00011_ clknet_leaf_25_clk_i memory\[40\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12264_ memory\[30\]\[10\] memory\[31\]\[10\] _06193_ _06470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_43_1200 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_120_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13251__S1 _02171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_32_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_107_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08958__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14003_ _01042_ clknet_leaf_164_clk_i memory\[59\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_147_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11215_ _05534_ _00627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_31_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1244 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12195_ _06401_ _06402_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_107_1289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput50 net50 data_o[19] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__10765__I0 _05016_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07176__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput61 net61 data_o[29] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__09592__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07630__I0 _03135_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11146_ _03359_ memory\[58\]\[24\] _05493_ _05498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_404_clk_i clknet_5_3__leaf_clk_i clknet_leaf_404_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_297_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11077_ _05461_ _00562_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12810__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10517__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09383__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10028_ _04629_ memory\[42\]\[26\] _04883_ _04890_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14905_ _01944_ clknet_leaf_70_clk_i memory\[35\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_160_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_601 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_14836_ _01875_ clknet_leaf_76_clk_i memory\[33\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11890__A1 _05699_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_176_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09135__I0 _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_419_clk_i clknet_5_2__leaf_clk_i clknet_leaf_419_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__07840__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_689 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11870__B _05687_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14767_ _01806_ clknet_leaf_128_clk_i memory\[31\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_175_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11979_ _05748_ _06183_ _06185_ _06188_ _06189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_15_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_85_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13718_ _03090_ _00776_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_156_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14698_ _01737_ clknet_leaf_169_clk_i memory\[2\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_74_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_907 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_85_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13649_ memory\[14\]\[31\] memory\[15\]\[31\] _05773_ _03036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_160_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_183_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07170_ _03118_ _03265_ _03306_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XANTENNA__08671__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_171_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_143_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_42_724 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_578 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_41_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15319_ _00278_ clknet_leaf_266_clk_i memory\[48\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_140_910 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_14_448 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_136_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_140_943 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_854 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_100_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09811_ _04774_ _02063_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_10_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_94_31 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_185_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10441__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09742_ _04737_ _02031_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06954_ net13 _03171_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_158_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_1240 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_09673_ _04616_ memory\[37\]\[20\] _04700_ _04701_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06885_ net3 _03117_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__13752__S _03074_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08624_ _04115_ _01535_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_55_1126 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__11881__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07750__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_46_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_77_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_89_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08555_ _04078_ _01503_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_178_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13622__A2 _02979_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_59_Left_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_49_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07688__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07506_ _03492_ _03504_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11633__A1 _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_542 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08486_ _03760_ memory\[21\]\[4\] _04037_ _04042_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_42_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_350 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_18_732 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_42_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07437_ memory\[49\]\[10\] _03329_ _03466_ _03467_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_130_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_21_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_383 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13386__A1 _05715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09677__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08581__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_545 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_31_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_190_865 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07368_ _03428_ _00966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_134_258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13199__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09107_ _04235_ memory\[2\]\[25\] _04380_ _04386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_72_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07299_ memory\[11\]\[11\] _03332_ _03390_ _03392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10995__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_60_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_103_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_115_483 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_111 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09038_ _04349_ _01715_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_14_993 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13233__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12116__B _05757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_68_Left_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_13_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12831__S _06751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10747__I0 _05066_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07925__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11000_ _05420_ _00526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11447__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_176_1221 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_142_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output51_I net51 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_201 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_142_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_19_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11547__S1 _05762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12951_ memory\[44\]\[20\] memory\[45\]\[20\] _02210_ _02349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11172__I0 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_172_1129 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__13662__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11902_ memory\[40\]\[5\] memory\[41\]\[5\] memory\[42\]\[5\] memory\[43\]\[5\] _05761_
+ _05762_ _06113_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_169_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15670_ _00629_ clknet_leaf_142_clk_i memory\[5\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11872__A1 _05690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_390_clk_i clknet_5_3__leaf_clk_i clknet_leaf_390_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_73_1226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12882_ memory\[40\]\[19\] memory\[41\]\[19\] memory\[42\]\[19\] memory\[43\]\[19\]
+ _06875_ _02217_ _02281_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XTAP_TAPCELL_ROW_29_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09117__I0 _04245_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_73_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_EDGE_ROW_77_Left_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14621_ _01660_ clknet_leaf_406_clk_i memory\[27\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11833_ memory\[44\]\[4\] memory\[45\]\[4\] _05749_ _06045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_96_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11182__S _05507_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_520 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14552_ _01591_ clknet_leaf_84_clk_i memory\[24\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11624__A1 _05741_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_67_153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11764_ memory\[40\]\[3\] memory\[41\]\[3\] memory\[42\]\[3\] memory\[43\]\[3\] _05761_
+ _05762_ _05977_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XPHY_EDGE_ROW_161_Right_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_55_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_82_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13503_ memory\[56\]\[29\] memory\[57\]\[29\] memory\[58\]\[29\] memory\[59\]\[29\]
+ _05711_ _03748_ _02892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_138_575 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_715 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10715_ _05269_ _00392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_181_810 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14483_ _01522_ clknet_leaf_105_clk_i memory\[22\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11695_ _05753_ _05908_ _05757_ _05909_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_55_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_181_832 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_597 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13434_ _02824_ net59 _02382_ _02825_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10646_ memory\[51\]\[13\] _03165_ _05229_ _05233_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_181_876 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_63_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13365_ _02371_ _02756_ _02373_ _02757_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__10526__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12805__I _05669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10577_ _05033_ memory\[50\]\[13\] _05192_ _05196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15104_ _00063_ clknet_leaf_439_clk_i memory\[42\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XPHY_EDGE_ROW_86_Left_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12316_ _06024_ _06516_ _06518_ _06520_ _06521_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__07851__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13296_ memory\[24\]\[25\] memory\[25\]\[25\] memory\[26\]\[25\] memory\[27\]\[25\]
+ _02363_ _02502_ _02689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12026__B _05722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_122_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_114_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15035_ _02074_ clknet_leaf_395_clk_i memory\[3\]\[31\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_107_1064 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_114_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12247_ _05667_ _06453_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07603__I0 _03197_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_343_clk_i clknet_5_8__leaf_clk_i clknet_leaf_343_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_12178_ _05732_ _06380_ _06382_ _06384_ _06385_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_120_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11357__S _05602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11129_ _03342_ memory\[58\]\[16\] _05482_ _05489_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09356__I0 _04212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_120_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_64_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_358_clk_i clknet_5_2__leaf_clk_i clknet_leaf_358_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__11863__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_976 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_149_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_91_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_154_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14819_ _01858_ clknet_leaf_402_clk_i memory\[33\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_626 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_148_317 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15799_ _00758_ clknet_leaf_59_clk_i net59 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_59_654 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11092__S _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_8_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_50_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08340_ net75 _03528_ _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XTAP_TAPCELL_ROW_177_3773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_175_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_177_3784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_47_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_698 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_15_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_131_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_564 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08271_ _03927_ _01370_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_15_1187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13368__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07222_ _03174_ _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_116_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_27_595 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07153_ _03203_ memory\[13\]\[25\] _03290_ _03296_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_375 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08095__I0 _03779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13320__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_70_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07084_ _03206_ memory\[16\]\[26\] _03251_ _03258_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_124_291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07842__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_930 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_125_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10729__I0 _05047_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_59_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_121_1028 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_1125 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_61_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_61_1196 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11267__S _05554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_81 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_96_1215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_35_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_35_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07986_ _03143_ _03764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XANTENNA_clkbuf_leaf_20_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09960__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12726__S0 _06582_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09725_ _04728_ _02023_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_06937_ _03158_ _00805_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11154__I0 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11854__A1 _05794_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_1081 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09656_ _04600_ memory\[37\]\[12\] _04689_ _04692_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07480__S _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_96_226 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08607_ _04105_ _01528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_26_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09587_ _04655_ _01958_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_136_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08538_ _03812_ memory\[21\]\[29\] _04059_ _04069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_245_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08469_ _04032_ _01463_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_9_261 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11730__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10500_ _05024_ memory\[4\]\[9\] _05145_ _05155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_108_759 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_135_556 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11480_ _05690_ _05695_ _05696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_33_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_98_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_98_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10431_ _05118_ _00259_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08086__I0 _03770_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10346__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10968__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09822__I1 _03205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_61_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_576 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_59_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13150_ _02319_ _02537_ _02544_ _02545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_59_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10362_ _05022_ memory\[47\]\[8\] _05073_ _05082_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_965 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_20_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_108_1351 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13657__S _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12101_ _05699_ _06299_ _06308_ _06309_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_TAPCELL_ROW_76_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12561__S _06557_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13081_ _02319_ _02468_ _02476_ _02477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_TAPCELL_ROW_76_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10293_ _05037_ memory\[46\]\[15\] _05027_ _05038_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_103_486 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07655__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09586__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12032_ _06240_ _06241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_0_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_109_18 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_72_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10081__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_206 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13983_ _01022_ clknet_leaf_329_clk_i memory\[59\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_176_1084 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15722_ _00681_ clknet_leaf_237_clk_i memory\[61\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12934_ memory\[8\]\[20\] memory\[9\]\[20\] memory\[10\]\[20\] memory\[11\]\[20\]
+ _06582_ _06721_ _02332_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__08486__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_125_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_16_Right_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__07390__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_150_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15653_ _00612_ clknet_leaf_312_clk_i memory\[5\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12865_ memory\[14\]\[19\] memory\[15\]\[19\] _02193_ _02264_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_34_1029 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__11704__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1344 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14604_ _01643_ clknet_leaf_124_clk_i memory\[26\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13598__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_68_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_157_136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11816_ _05681_ _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15584_ _00543_ clknet_leaf_324_clk_i memory\[57\]\[4\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_51_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12796_ _06717_ _02194_ _02195_ _02196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_141_16 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09510__I0 _04606_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_173_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14535_ _01574_ clknet_leaf_175_clk_i memory\[24\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_56_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11747_ memory\[14\]\[3\] memory\[15\]\[3\] _05720_ _05960_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_155_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_126_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_155_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_148_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14466_ _01505_ clknet_leaf_357_clk_i memory\[22\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_12_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_342 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11678_ _05719_ _05891_ _05722_ _05892_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_172_3681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_116_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_172_3692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12022__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13417_ _02336_ _02800_ _02807_ _02808_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_181_684 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10629_ memory\[51\]\[5\] _03140_ _05218_ _05224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11456__S0 _05670_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10256__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_109_1115 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_180_172 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_25_Right_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_14397_ _01436_ clknet_leaf_358_clk_i memory\[20\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_144_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_52_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_133_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07824__I0 _03221_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13348_ _02739_ _02740_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
Xclkbuf_leaf_282_clk_i clknet_5_12__leaf_clk_i clknet_leaf_282_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_45_1169 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13279_ memory\[38\]\[25\] memory\[39\]\[25\] _05662_ _02672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07565__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15018_ _02057_ clknet_leaf_249_clk_i memory\[3\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_122_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09577__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11595__B _05807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12956__S0 _06875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12270__I _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07840_ _03144_ memory\[7\]\[6\] _03675_ _03682_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07364__I _03414_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09329__I0 _04185_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09780__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_75_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_297_clk_i clknet_5_15__leaf_clk_i clknet_leaf_297_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA_clkbuf_leaf_194_clk_i_I clknet_5_31__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07771_ _03645_ _01152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XPHY_EDGE_ROW_34_Right_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_09510_ _04606_ memory\[35\]\[15\] _04596_ _04607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_179_3813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_95_1270 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__08396__S _03987_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11836__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_179_3824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_32 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_09441_ _04229_ memory\[34\]\[22\] _04560_ _04563_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xclkbuf_leaf_220_clk_i clknet_5_27__leaf_clk_i clknet_leaf_220_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_8_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_91_1178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13589__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09372_ _04526_ _01872_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_192_905 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_19_315 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09257__A2 _03305_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_46_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__09501__I0 _04600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08323_ _03955_ _01394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_46_123 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12646__S _06845_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_117_512 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_7_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_523 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12800__A3 _02199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08254_ _03800_ memory\[17\]\[23\] _03915_ _03919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_61_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_235_clk_i clknet_5_15__leaf_clk_i clknet_leaf_235_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_1231 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_43_Right_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09020__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_27_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_7_787 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07205_ memory\[39\]\[10\] _03329_ _03330_ _03331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_132_515 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12013__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08068__I0 _03746_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10166__S _04955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08185_ _03882_ _01329_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_537 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07136_ _03178_ memory\[13\]\[17\] _03279_ _03287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_43_896 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_113_762 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07067_ _03181_ memory\[16\]\[18\] _03240_ _03249_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_37_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_37_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_140_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_11_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13513__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_101_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_54_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11375__I0 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_10_281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_EDGE_ROW_52_Right_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_177_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07969_ _03746_ memory\[12\]\[0\] _03752_ _03753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__11127__I0 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11725__S _05868_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09708_ _04719_ _02015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_10980_ _05398_ _05410_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_74_1354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09639_ _04583_ memory\[37\]\[4\] _04678_ _04683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_35_1338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_66_911 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12650_ _06848_ _06849_ _06707_ _06850_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_TAPCELL_ROW_137_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11601_ _05690_ _05815_ _05816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_65_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_396_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_66_966 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12581_ _06155_ _06776_ _06778_ _06781_ _06782_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_148_681 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_61_Right_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_81_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_92_251 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14320_ _01359_ clknet_leaf_115_clk_i memory\[17\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_318 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11532_ _05747_ _05748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_68_1114 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_178 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_68_1136 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_11_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_78_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14251_ _01290_ clknet_leaf_198_clk_i memory\[15\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12004__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_162_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_11463_ memory\[52\]\[0\] memory\[53\]\[0\] _05678_ _05679_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_80_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_145_1326 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13202_ _06848_ _02595_ _05791_ _02596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_34_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09865__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07806__I0 _03194_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12555__A2 _06748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_150_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_345 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_145_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10414_ _05004_ memory\[48\]\[0\] _05109_ _05110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14182_ _01221_ clknet_leaf_205_clk_i memory\[19\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11394_ _03334_ memory\[62\]\[12\] _05627_ _05630_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_21_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_74_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_389 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13133_ _06838_ _02527_ _02528_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_10345_ _05072_ _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__07282__I1 _03315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_104_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_111_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_111_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_143_1072 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09559__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13504__A1 _05710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_103_294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13064_ _06831_ _02455_ _02457_ _02459_ _02460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_10276_ _03155_ _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_104_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_44_1191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_70_Right_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_12015_ _05651_ _06216_ _06223_ _06224_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__08231__I0 _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_79_1243 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11818__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13966_ _01005_ clknet_leaf_258_clk_i memory\[49\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_109_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_177_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09105__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_186_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15705_ _00664_ clknet_leaf_382_clk_i memory\[60\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12917_ memory\[48\]\[20\] memory\[49\]\[20\] memory\[50\]\[20\] memory\[51\]\[20\]
+ _06699_ _06839_ _02315_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__12491__A1 _06279_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13897_ _00936_ clknet_leaf_212_clk_i memory\[11\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_157_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_17_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_88_579 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_1130 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_69_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_75_207 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_115_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_968 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_152_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15636_ _00595_ clknet_leaf_166_clk_i memory\[58\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_69_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12848_ memory\[52\]\[19\] memory\[53\]\[19\] _06832_ _02247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08944__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_28_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_174_3721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_173_404 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_8_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__13666__S1 _05694_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_115_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_51_1151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_150_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15567_ _00526_ clknet_leaf_243_clk_i memory\[56\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_167_990 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12779_ _06835_ _02177_ _02178_ _02179_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_185_1106 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_185_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14518_ _01557_ clknet_leaf_91_clk_i memory\[23\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_126_331 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15498_ _00457_ clknet_leaf_239_clk_i memory\[54\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_25_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_117_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_4_713 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14449_ _01488_ clknet_leaf_99_clk_i memory\[21\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_181_481 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_25_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_3_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_52_660 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_101_41 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_12_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08470__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09990_ _04591_ memory\[42\]\[8\] _04861_ _04870_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10714__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08941_ _04298_ _01669_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_86_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_0_985 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08222__I0 _03768_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08872_ _04203_ memory\[26\]\[10\] _04261_ _04262_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_32_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09970__I0 _04639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07823_ _03672_ _01177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_5_15__f_clk_i clknet_2_1_0_clk_i clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07754_ _03218_ memory\[63\]\[30\] _03602_ _03636_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08918__I _04285_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09722__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_189_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__12482__A1 _06639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07685_ _03599_ _01112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_09424_ _04212_ memory\[34\]\[14\] _04549_ _04554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_456 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_192_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_177_776 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_165_927 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_730 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_489 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_165_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12234__A1 _06028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09355_ _04517_ _01864_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_191_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_174_clk_i clknet_5_28__leaf_clk_i clknet_leaf_174_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__12376__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11280__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_48_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_75_774 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08306_ _03946_ _01386_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10096__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_129_191 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09286_ _04210_ memory\[32\]\[13\] _04477_ _04481_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_7_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08237_ _03783_ memory\[17\]\[15\] _03904_ _03910_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_95_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_132_312 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_334 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_43_671 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09685__S _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_559 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_189_clk_i clknet_5_29__leaf_clk_i clknet_leaf_189_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_166_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08168_ _03873_ _01321_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10548__A1 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_30_321 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_120_518 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__07413__A1 _03451_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07119_ _03153_ memory\[13\]\[9\] _03268_ _03278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_570 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_120_529 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08099_ _03783_ memory\[15\]\[15\] _03830_ _03836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_113_581 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_24_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09484__I _03146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_899 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10130_ _04932_ _04944_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_101_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_30_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_112_clk_i clknet_5_23__leaf_clk_i clknet_leaf_112_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_100_264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10061_ _04907_ _00100_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07933__S _03722_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10020__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13820_ _00859_ clknet_leaf_373_clk_i memory\[13\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_127_clk_i clknet_5_29__leaf_clk_i clknet_leaf_127_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_98_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08828__I _03202_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_187_507 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_3_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09713__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13751_ _03107_ _00792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_1027 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_721 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12473__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10963_ _05401_ _00508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_39_1282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_98_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__13670__S _02495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_167_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12702_ memory\[62\]\[17\] memory\[63\]\[17\] _06557_ _02103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08764__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13682_ _05760_ _03068_ _03069_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_57_229 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_67_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_183_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10894_ memory\[55\]\[1\] _03128_ _05363_ _05365_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_104_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15421_ _00380_ clknet_leaf_345_clk_i memory\[52\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_191_4054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_168_798 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12633_ memory\[52\]\[16\] memory\[53\]\[16\] _06832_ _06833_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_752 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12286__S _06491_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_54_914 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_152_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15352_ _00311_ clknet_leaf_44_clk_i memory\[4\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_152_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_54_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12564_ _06279_ _06764_ _06765_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_142_clk_i_I clknet_5_19__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14303_ _01342_ clknet_leaf_350_clk_i memory\[17\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_301 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11515_ _03304_ _05731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_0_1155 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15283_ _00242_ clknet_leaf_40_clk_i memory\[47\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_145_1101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12495_ memory\[54\]\[14\] memory\[55\]\[14\] _06421_ _06697_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_151_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_0_1166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07179__I _03131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_14234_ _01273_ clknet_leaf_30_clk_i memory\[12\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11446_ _05661_ _05662_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_123_367 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08452__I0 _03793_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14165_ _01204_ clknet_leaf_136_clk_i memory\[7\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_215 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12813__I _05681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10534__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11377_ _03317_ memory\[62\]\[4\] _05616_ _05621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_104_592 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09394__I _04537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13116_ _02367_ _02507_ _02509_ _02511_ _02512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_81_1188 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10328_ _05061_ _00213_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14096_ _01135_ clknet_leaf_133_clk_i memory\[63\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12034__B _06177_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_13_Left_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_167_3591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13047_ _02398_ _02413_ _02428_ _02443_ _02444_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__12387__S1 _06454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10259_ _05014_ memory\[46\]\[4\] _05006_ _05015_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10011__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09952__I0 _04621_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_128_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11365__S _05579_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13336__S0 _02473_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_67_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14998_ _02037_ clknet_leaf_66_clk_i memory\[38\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_710 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_57_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12464__A1 _06325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13949_ _00988_ clknet_leaf_345_clk_i memory\[49\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_72_56 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_754 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_91_clk_i clknet_5_20__leaf_clk_i clknet_leaf_91_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_48_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_5_8__f_clk_i_I clknet_2_1_0_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07470_ memory\[49\]\[26\] _03363_ _03477_ _03484_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_147_916 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_607 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_EDGE_ROW_22_Left_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_5_1022 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_432 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_629 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_147_949 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_146_426 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15619_ _00578_ clknet_leaf_321_clk_i memory\[58\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_9_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12196__S _06062_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_173_212 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_286 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_158_297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09140_ _04403_ _01763_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_29_487 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12209__B _06001_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_44_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09071_ _04199_ memory\[2\]\[8\] _04358_ _04367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_115_835 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07494__I1 _03317_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08691__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_47_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08022_ _03788_ _01260_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_71_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_868 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_141_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_12_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08443__I0 _03785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_187_3967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_31_Left_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_90_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10250__I0 _05008_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_86 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_25_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_12_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_344_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09973_ _04860_ _04861_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_08924_ _04289_ _01661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__13495__A3 _02884_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_44_clk_i clknet_5_18__leaf_clk_i clknet_leaf_44_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__09943__I0 _04612_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08855_ _04187_ memory\[26\]\[2\] _04250_ _04253_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_98_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07806_ _03194_ memory\[6\]\[22\] _03661_ _03664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_2_Right_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_08786_ _04206_ memory\[25\]\[11\] _04204_ _04207_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_88_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input13_I data_i[15] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_88_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07737_ _03627_ _01136_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12455__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_59_clk_i clknet_5_17__leaf_clk_i clknet_leaf_59_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XPHY_EDGE_ROW_40_Left_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_TAPCELL_ROW_49_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13490__S _05754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1324 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07668_ _03191_ memory\[10\]\[21\] _03589_ _03591_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_165_702 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09407_ _04195_ memory\[34\]\[6\] _04538_ _04545_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10619__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07599_ _03191_ memory\[0\]\[21\] _03552_ _03554_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_137_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10069__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_1190 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__08383__I _03964_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09338_ _04508_ _01856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_164_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1145 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_871 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_62_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_164_289 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_35_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_117_161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09269_ _04193_ memory\[32\]\[5\] _04466_ _04472_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_69_1264 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_22_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_11300_ _05579_ _05580_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_12280_ memory\[16\]\[10\] memory\[17\]\[10\] memory\[18\]\[10\] memory\[19\]\[10\]
+ _06342_ _06485_ _06486_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_161_996 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_105_378 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_181_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11231_ _05542_ _05543_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__10354__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11162_ _03266_ _03528_ _05506_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
X_10113_ _04935_ _00124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_8_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_8_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__13566__S0 _05711_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11093_ _05469_ _00570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07663__S _03578_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10044_ _04577_ memory\[43\]\[1\] _04897_ _04899_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14921_ _01960_ clknet_leaf_36_clk_i memory\[36\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_145_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11185__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14852_ _01891_ clknet_leaf_400_clk_i memory\[34\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_69_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13803_ _00842_ clknet_leaf_206_clk_i memory\[16\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_193_4105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14783_ _01822_ clknet_leaf_420_clk_i memory\[32\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11995_ _05794_ _06204_ _06205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_123_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11913__S _05785_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13734_ _03353_ memory\[9\]\[21\] _03097_ _03099_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_58_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08494__S _04037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10946_ memory\[55\]\[26\] _03205_ _05385_ _05392_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_42_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_13665_ _05682_ _03051_ _05722_ _03052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__13413__B _02352_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_128_437 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10877_ _05060_ memory\[54\]\[26\] _05348_ _05355_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_54_700 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12616_ memory\[16\]\[15\] memory\[17\]\[15\] memory\[18\]\[15\] memory\[19\]\[15\]
+ _06342_ _06485_ _06817_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_156_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15404_ _00363_ clknet_leaf_258_clk_i memory\[51\]\[16\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_155_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_1252 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13596_ memory\[32\]\[30\] memory\[33\]\[30\] memory\[34\]\[30\] memory\[35\]\[30\]
+ _05670_ _05671_ _02984_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA_clkbuf_leaf_293_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_15335_ _00294_ clknet_leaf_242_clk_i memory\[4\]\[11\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12547_ memory\[20\]\[14\] memory\[21\]\[14\] _06477_ _06749_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07476__I1 _03369_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_941 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07838__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15266_ _00225_ clknet_leaf_404_clk_i memory\[47\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_83_1228 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12478_ memory\[16\]\[13\] memory\[17\]\[13\] memory\[18\]\[13\] memory\[19\]\[13\]
+ _06342_ _06485_ _06681_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XANTENNA__12057__S0 _05795_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_169_3620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14217_ _01256_ clknet_leaf_217_clk_i memory\[12\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_123_175 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_22_641 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11429_ _03369_ memory\[62\]\[29\] _05638_ _05648_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_15197_ _00156_ clknet_leaf_436_clk_i memory\[45\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_6_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__10232__I0 _04629_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1_568 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14148_ _01187_ clknet_leaf_286_clk_i memory\[7\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_67_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_123_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_69 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06970_ net17 _03183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_14079_ _01118_ clknet_leaf_310_clk_i memory\[63\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08669__S _04132_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_184_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_input5_I address_i[4] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07573__S _03530_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_182_3875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12685__A1 _06607_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_158_1347 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_20_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_119_1309 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08640_ memory\[23\]\[12\] _03334_ _04121_ _04124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_179_805 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_EDGE_ROW_175_Right_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12780__S1 _06839_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_816 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08571_ _03777_ memory\[22\]\[12\] _04084_ _04087_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_53_1010 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10299__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_178_359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_07522_ _03512_ _01036_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_18_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_159_562 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_07453_ memory\[49\]\[18\] _03346_ _03466_ _03475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_174_521 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10439__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__06911__I0 _03138_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_779 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07384_ _03436_ _00974_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_123_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_18_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_44_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_587 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09123_ _04181_ memory\[30\]\[0\] _04394_ _04395_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_621 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_115_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07748__S _03625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_40_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_09054_ _04357_ _04358_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_89_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_1140 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11778__B _05792_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_142_462 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_60_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08005_ _03162_ _03777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_103_838 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08416__I0 _03758_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10174__S _04932_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_130_646 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_1281 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_64_1161 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_163_1097 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_679 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_5_30__f_clk_i clknet_2_3_0_clk_i clknet_5_30__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_12_195 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11069__I _05434_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_102_1313 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13548__S0 _02363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10902__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09956_ _04625_ memory\[41\]\[24\] _04847_ _04852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_110_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08579__S _04084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_5_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_99_1257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_1357 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08907_ _04239_ memory\[26\]\[27\] _04272_ _04280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09916__I0 _04585_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09887_ _04815_ _00018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08838_ _04241_ memory\[25\]\[28\] _04225_ _04242_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_142_Right_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__12428__A1 _06272_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08769_ _03143_ _04195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__12829__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_140_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_71_1110 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10800_ _05314_ _00432_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_140_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_68_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11780_ _05794_ _05992_ _05993_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__07155__I0 _03206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_184_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09203__S _04430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_64_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_101_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_806 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10731_ _05050_ memory\[52\]\[21\] _05276_ _05278_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_193_830 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177_381 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11532__I _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_81_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_165_554 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_76_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_81_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13450_ _02302_ _02832_ _02839_ _02840_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
X_10662_ _05241_ _00367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_960 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_119_982 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12401_ memory\[28\]\[12\] memory\[29\]\[12\] _06604_ _06605_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_766 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_15_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12600__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13381_ _02771_ _02772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__07458__I1 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_106_632 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10593_ _05204_ _00335_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_35_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15120_ _00079_ clknet_leaf_8_clk_i memory\[42\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12332_ _06445_ _06529_ _06536_ _06537_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__10462__I0 _05054_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_105_142 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_51_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15051_ _00010_ clknet_leaf_33_clk_i memory\[40\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13156__A2 _02550_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12263_ _06468_ _06469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__10084__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12203__I1 net71 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_181_1186 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_14002_ _01041_ clknet_leaf_163_clk_i memory\[59\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07457__I _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11214_ _03359_ memory\[5\]\[24\] _05529_ _05534_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09873__S _04800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_147_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_82_1283 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__09080__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12194_ memory\[20\]\[9\] memory\[21\]\[9\] _05785_ _06401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_147_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xoutput40 net40 data_o[0] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XFILLER_0_43_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13395__S _05769_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput51 net51 data_o[1] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__11908__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput62 net62 data_o[2] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
X_11145_ _05497_ _00594_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09672__I _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_179_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_11076_ _05054_ memory\[57\]\[23\] _05457_ _05461_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12667__A1 _06450_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_125_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11707__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10027_ _04889_ _00084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14904_ _01943_ clknet_leaf_70_clk_i memory\[35\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07394__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_160_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12419__A1 _06570_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14835_ _01874_ clknet_leaf_75_clk_i memory\[33\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12739__S _06596_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_121_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_188_657 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_37_1049 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_121_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11643__S _05789_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14766_ _01805_ clknet_leaf_127_clk_i memory\[31\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_153_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_11978_ _05760_ _06187_ _06188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__09113__S _04380_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13717_ _03336_ memory\[9\]\[13\] _03086_ _03090_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_86_677 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10929_ memory\[55\]\[18\] _03180_ _05374_ _05383_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14697_ _01736_ clknet_leaf_169_clk_i memory\[2\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10259__S _05006_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_128_234 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_176 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_768 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_128_256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_73_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08952__S _04297_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13648_ _03034_ _03035_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__07449__I1 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12474__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_703 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13579_ memory\[6\]\[30\] memory\[7\]\[30\] _05795_ _02967_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_492 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_125_963 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10453__I0 _05045_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08751__I _04182_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15318_ _00277_ clknet_leaf_267_clk_i memory\[48\]\[26\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_124_451 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_2_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_48_1167 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15249_ _00208_ clknet_leaf_43_clk_i memory\[46\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_1_332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10205__I0 _04602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_184_3915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_99_Right_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_140_999 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09071__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_156 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09810_ memory\[3\]\[20\] _03186_ _04773_ _04774_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_10_655 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10722__S _05265_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09741_ _04616_ memory\[38\]\[20\] _04736_ _04737_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06953_ _03170_ _00809_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12658__A1 _06717_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_87 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09672_ _04677_ _04700_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_94_1121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_06884_ net2 _03116_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XFILLER_0_94_1143 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_1154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_97_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_178_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08623_ memory\[23\]\[4\] _03317_ _04110_ _04115_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_1116 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_85_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__12649__S _06431_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08554_ _03760_ memory\[22\]\[4\] _04073_ _04078_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_166_307 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_46_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_193_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_166_329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07505_ _03503_ _01028_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_187_690 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08485_ _04041_ _01470_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_65_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_42_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__09958__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_76_187 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07436_ _03454_ _03466_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_64_338 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_21_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_80_809 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_169_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_21_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_73_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_45_552 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07367_ _03160_ memory\[8\]\[11\] _03426_ _03428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_872 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_189_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09106_ _04385_ _01747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_17_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07478__S _03454_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_760 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_60_533 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07298_ _03391_ _00933_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_33_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09037_ _04233_ memory\[28\]\[24\] _04344_ _04349_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_102_101 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_66_1278 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_102_134 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_131_977 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09693__S _04677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12441__S0 _06020_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_57_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_241_clk_i_I clknet_5_13__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_141_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09939_ _04608_ memory\[41\]\[16\] _04836_ _04843_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_142_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11527__I _03747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_142_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12950_ _02337_ _02340_ _02343_ _02347_ _02348_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA_output44_I net44 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_137_1239 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11901_ _05753_ _06111_ _05757_ _06112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_12881_ _02213_ _02279_ _06461_ _02280_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12559__S _06273_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11463__S _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_29_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_29_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11832_ _05732_ _06038_ _06041_ _06043_ _06044_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
X_14620_ _01659_ clknet_leaf_390_clk_i memory\[27\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07128__I0 _03166_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_185_627 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_138_510 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14551_ _01590_ clknet_leaf_80_clk_i memory\[24\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_36_1071 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_96_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08876__I0 _04208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11763_ _05753_ _05975_ _05757_ _05976_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__10079__S _04908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12821__A1 _06445_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10714_ _05033_ memory\[52\]\[13\] _05265_ _05269_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_13502_ _05705_ _02890_ _05756_ _02891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_14482_ _01521_ clknet_leaf_101_clk_i memory\[22\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_166_874 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_166_885 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11694_ memory\[46\]\[2\] memory\[47\]\[2\] _05907_ _05908_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_55_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_126_727 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_1356 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_193_682 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_13433_ _02778_ _02793_ _02808_ _02823_ _02824_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_0_10_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10645_ _05232_ _00359_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_119_790 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10807__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07388__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_24_725 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_51_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10435__I0 _05026_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13364_ memory\[22\]\[26\] memory\[23\]\[26\] _05754_ _02756_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_109_1319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10576_ _05195_ _00327_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_180_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_2_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_134_782 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12315_ _06031_ _06519_ _06520_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_15103_ _00062_ clknet_leaf_439_clk_i memory\[42\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_23_268 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_122_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13295_ _02498_ _02687_ _02086_ _02688_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_45_1329 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15034_ _02073_ clknet_leaf_28_clk_i memory\[3\]\[30\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_114_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12246_ _06450_ _06451_ _06177_ _06452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XTAP_TAPCELL_ROW_114_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_43_1042 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12177_ _05741_ _06383_ _06384_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__10542__S _05167_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_20_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_177_1019 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11560__A1 _05772_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11128_ _05488_ _00586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08012__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10341__I _03220_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11059_ _05037_ memory\[57\]\[15\] _05446_ _05452_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07367__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_79_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07851__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12469__S _06193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_188_443 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10910__I1 _03152_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11373__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_99_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_8_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_188_465 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13065__A1 _02302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14818_ _01857_ clknet_leaf_429_clk_i memory\[33\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA_clkbuf_leaf_443_clk_i_I clknet_5_1__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07119__I0 _03153_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15798_ _00757_ clknet_leaf_58_clk_i net58 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_118_1183 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_188_498 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_147_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_114_1036 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_87_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_177_3774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08867__I0 _04199_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14749_ _01788_ clknet_leaf_391_clk_i memory\[31\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_46_305 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_191_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_177_3785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_157_863 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09778__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08270_ _03816_ memory\[17\]\[31\] _03892_ _03927_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_73_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_190_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_362 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_6_402 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_129_598 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_13_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_89_1256 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07221_ _03341_ _00906_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_144_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_15_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_117_749 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_190_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_6_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_55_894 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_172_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__10426__I0 _05018_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07152_ _03295_ _00883_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09292__I0 _04216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_131_218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_769 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13099__I _05655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12217__B _06287_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_65 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_30_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_14_257 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07083_ _03257_ _00852_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12932__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_160_1012 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_23_780 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_113_988 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_11_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_39_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_26_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_100_649 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_10_463 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09018__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_22_1159 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_35_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07985_ _03763_ _01248_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_96_1227 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09724_ _04600_ memory\[38\]\[12\] _04725_ _04728_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12726__S1 _06721_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_06936_ _03156_ memory\[14\]\[10\] _03157_ _03158_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__08857__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07358__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09655_ _04691_ _01990_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08606_ _03812_ memory\[22\]\[29\] _04095_ _04105_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_171_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_167_605 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_26_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08656__I _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13056__A1 _02170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_26_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_78_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09586_ _04598_ memory\[36\]\[11\] _04653_ _04655_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_78_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_171_1185 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08537_ _04068_ _01495_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_49_165 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_400 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72_1293 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_64_113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08592__S _04095_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08468_ _03810_ memory\[20\]\[28\] _04023_ _04032_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_163_822 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_174_170 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07419_ _03457_ _00988_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_52_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08399_ _03995_ _01430_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_403_clk_i clknet_5_2__leaf_clk_i clknet_leaf_403_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__10627__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_354 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09487__I _03149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10430_ _05022_ memory\[48\]\[8\] _05109_ _05118_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_98_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_61_842 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_98_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_6_980 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07001__S _03188_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_59_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11090__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_143_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10361_ _05081_ _00226_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_27_1015 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_104_944 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_59_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_1075 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11790__A1 _05660_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12100_ _06024_ _06301_ _06305_ _06307_ _06308_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_13080_ _06713_ _02470_ _02472_ _02475_ _02476_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__09035__I0 _04231_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_418_clk_i clknet_5_2__leaf_clk_i clknet_leaf_418_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_76_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_130_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10292_ _03171_ _05037_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_12031_ memory\[36\]\[7\] memory\[37\]\[7\] _05733_ _06240_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10362__S _05073_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07597__I0 _03187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_392_clk_i_I clknet_5_3__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11542__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13295__A1 _02498_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13982_ _01021_ clknet_leaf_326_clk_i memory\[59\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08767__S _04183_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15721_ _00680_ clknet_leaf_235_clk_i memory\[61\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12933_ _06717_ _02330_ _02195_ _02331_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_0_77_1182 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11193__S _05518_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_154_1361 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08566__I _04072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13047__A1 _02398_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15652_ _00611_ clknet_leaf_282_clk_i memory\[5\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12864_ _02262_ _02263_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_150_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_73_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_38_1199 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14603_ _01642_ clknet_leaf_185_clk_i memory\[26\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11815_ _06026_ _06027_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_12795_ _05664_ _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_15583_ _00542_ clknet_leaf_326_clk_i memory\[57\]\[3\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_29_839 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_83_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09598__S _04653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14534_ _01573_ clknet_leaf_175_clk_i memory\[24\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11746_ _05958_ _05959_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_172_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_155_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_50_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_55_146 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_155_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_138_384 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13421__B _05665_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14465_ _01504_ clknet_leaf_351_clk_i memory\[22\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11677_ memory\[14\]\[2\] memory\[15\]\[2\] _05720_ _05891_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12816__I _05689_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_165_192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_12_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_12_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_TAPCELL_ROW_172_3682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10408__I0 _05068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_116_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_180_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_172_3693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10628_ _05223_ _00351_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13416_ _02209_ _02802_ _02804_ _02806_ _02807_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XTAP_TAPCELL_ROW_116_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_153_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14396_ _01435_ clknet_leaf_361_clk_i memory\[20\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_84_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_183_1045 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11456__S1 _05671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_183_1056 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_49_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_133_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_45_1104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13347_ memory\[44\]\[26\] memory\[45\]\[26\] _02210_ _02739_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12752__S _06477_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_133_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10559_ _05186_ _00319_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_49_1284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12573__A3 _06773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_374 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_80_1006 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11781__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_1017 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_161_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__07846__S _03675_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09026__I0 _04222_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13278_ _02670_ _02671_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_110_936 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15017_ _02056_ clknet_leaf_249_clk_i memory\[3\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12229_ _06162_ _06434_ _06435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__12956__S1 _02217_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07588__I0 _03175_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_137_clk_i_I clknet_5_22__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07770_ _03141_ memory\[6\]\[5\] _03639_ _03645_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_159_1272 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__08677__S _04109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_179_3814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_56_1222 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_179_3825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_91_1113 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09440_ _04562_ _01904_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13038__A1 _06603_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_52_1108 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_56_1277 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_148_104 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07760__I0 _03111_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_91_66 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_75_901 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_47_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09371_ _04227_ memory\[33\]\[21\] _04524_ _04526_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_87_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_176_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_192_917 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_08322_ _03800_ memory\[18\]\[23\] _03951_ _03955_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_75_956 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_74_444 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09301__S _04488_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08253_ _03918_ _01361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_28_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_117_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10447__S _05120_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_166_1210 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_28_883 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_34_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_105_708 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_07204_ _03308_ _03330_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
X_08184_ _03798_ memory\[29\]\[22\] _03879_ _03882_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_131_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__09265__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_376 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_544 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1265 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_144_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_132_527 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_144_398 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_566 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07135_ _03286_ _00875_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11072__I0 _05050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10246__I _05005_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_15_599 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_71_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07756__S _03602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07066_ _03248_ _00844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_37_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_93_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11278__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_11_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__10182__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11524__A1 _05736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_54_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__10910__S _05363_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07968_ _03751_ _03752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_09707_ _04583_ memory\[38\]\[4\] _04714_ _04719_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_06919_ _03144_ memory\[14\]\[6\] _03126_ _03145_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_07899_ _03713_ _01212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_134_1209 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09638_ _04682_ _01982_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__13029__A1 _02216_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_547 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_179_262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_179_284 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_168_947 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09569_ _04581_ memory\[36\]\[3\] _04642_ _04646_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_66_923 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_155_608 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11600_ memory\[48\]\[1\] memory\[49\]\[1\] memory\[50\]\[1\] memory\[51\]\[1\] _05692_
+ _05694_ _05815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA_clkbuf_leaf_339_clk_i_I clknet_5_9__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_182_405 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_65_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_12580_ _06162_ _06780_ _06781_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_137_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_33_1052 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_38_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_182_427 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_342_clk_i clknet_5_8__leaf_clk_i clknet_leaf_342_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_93_764 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_108_524 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_11531_ _05652_ _05747_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_12
XFILLER_0_108_535 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_33_1096 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_263 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_343 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11540__I _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14250_ _01289_ clknet_leaf_201_clk_i memory\[15\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11462_ _05677_ _05678_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_68_1148 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_78_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_190_471 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_110_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_151_836 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13201_ memory\[6\]\[24\] memory\[7\]\[24\] _02322_ _02595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_33_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10413_ _05108_ _05109_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__11063__I0 _05041_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14181_ _01220_ clknet_leaf_368_clk_i memory\[19\]\[9\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_150_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11393_ _05629_ _00710_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_357_clk_i clknet_5_8__leaf_clk_i clknet_leaf_357_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_104_741 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_150_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11763__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07666__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13132_ memory\[48\]\[23\] memory\[49\]\[23\] memory\[50\]\[23\] memory\[51\]\[23\]
+ _06699_ _06839_ _02527_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__09008__I0 _04203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10344_ _03306_ _04787_ _05072_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_81_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_TAPCELL_ROW_111_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_108_1171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_103_273 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10092__S _04919_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13063_ _06838_ _02458_ _02459_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_40_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10275_ _05025_ _00196_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_12014_ _06142_ _06218_ _06220_ _06222_ _06223_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_104_1068 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_121_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13268__A1 _06844_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_40_1089 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_136_28 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__07990__I0 _03766_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13416__B _02804_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_88_503 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13965_ _01004_ clknet_leaf_257_clk_i memory\[49\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_109_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_159_903 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_15704_ _00663_ clknet_leaf_383_clk_i memory\[60\]\[28\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__10877__I0 _05060_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12916_ _06835_ _02313_ _02178_ _02314_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_13896_ _00935_ clknet_leaf_215_clk_i memory\[11\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07742__I0 _03200_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_157_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_150_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_17_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15635_ _00594_ clknet_leaf_164_clk_i memory\[58\]\[23\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_17_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_57_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12747__S _02084_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_614 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12847_ _02163_ _02241_ _02243_ _02245_ _02246_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_0_158_457 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_174_3722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_174_3733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_174_939 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15566_ _00525_ clknet_leaf_246_clk_i memory\[56\]\[18\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_5_1259 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09495__I0 _04595_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_57_978 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12778_ _05686_ _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_83_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_139_693 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_185_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14517_ _01556_ clknet_leaf_105_clk_i memory\[23\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11729_ _05654_ _05937_ _05939_ _05941_ _05942_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_15497_ _00456_ clknet_leaf_290_clk_i memory\[54\]\[13\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_182_961 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_154_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_182_994 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14448_ _01487_ clknet_leaf_100_clk_i memory\[21\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09247__I0 _04239_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_387 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_3_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12990__B _06690_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_63_clk_i_I clknet_5_16__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_80_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_142_869 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_141_346 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14379_ _01418_ clknet_leaf_200_clk_i memory\[1\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__07576__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10801__I0 _05052_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_51_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_0_920 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11098__S _05471_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08940_ _04203_ memory\[27\]\[10\] _04297_ _04298_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09791__S _04762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11357__I1 _03208_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_110_788 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08871_ _04249_ _04261_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_97_1311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_99 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_TAPCELL_ROW_32_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07822_ _03218_ memory\[6\]\[30\] _03638_ _03672_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_288_clk_i_I clknet_5_15__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13259__A1 _06838_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_58_1328 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_93_1208 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07981__I0 _03760_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07753_ _03635_ _01144_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08200__S _03856_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07684_ _03215_ memory\[10\]\[29\] _03589_ _03599_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_149_413 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12482__A2 _06654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_149_424 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09423_ _04553_ _01896_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_172_1291 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_165_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12657__S _06302_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_340_clk_i_I clknet_5_8__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_59_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_09354_ _04210_ memory\[33\]\[13\] _04513_ _04517_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13431__A1 _02367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08305_ _03783_ memory\[18\]\[15\] _03940_ _03946_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09031__S _04344_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10245__A1 _03124_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13061__B _02178_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09285_ _04480_ _01831_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11993__A1 _05788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08236_ _03909_ _01353_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__09966__S _04847_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_95_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_166_1051 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_127_1002 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_16_864 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13488__S _02368_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_144_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_15_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_08167_ _03781_ memory\[29\]\[14\] _03868_ _03873_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09789__I1 _03155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_31_812 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_166_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07486__S _03493_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_132_379 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_67_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07118_ _03277_ _00867_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_63_1034 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08098_ _03835_ _01289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__12405__B _06195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_EDGE_ROW_189_Right_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_101_744 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_07049_ _03239_ _00836_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_41_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_10060_ _04593_ memory\[43\]\[9\] _04897_ _04907_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12170__A1 _06024_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10640__S _05229_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07972__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1120 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__08110__S _03841_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_138_1153 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_3_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_3_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13750_ _03369_ memory\[9\]\[29\] _03097_ _03107_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_10962_ _05008_ memory\[56\]\[1\] _05399_ _05401_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_97_333 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_1294 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_12701_ _02101_ _02102_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_0_39_912 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_906 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10893_ _05364_ _00475_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_13681_ memory\[16\]\[31\] memory\[17\]\[31\] memory\[18\]\[31\] memory\[19\]\[31\]
+ _05761_ _05762_ _03068_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_38_411 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_281_clk_i clknet_5_12__leaf_clk_i clknet_leaf_281_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_104_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15420_ _00379_ clknet_leaf_332_clk_i memory\[52\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_38_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_104_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_191_4055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_12632_ _05677_ _06832_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_112_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11284__I0 _03361_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_152_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_66_786 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12563_ memory\[56\]\[15\] memory\[57\]\[15\] memory\[58\]\[15\] memory\[59\]\[15\]
+ _06138_ _06280_ _06764_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
X_15351_ _00310_ clknet_leaf_150_clk_i memory\[4\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_0_1112 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_109_877 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14302_ _01341_ clknet_leaf_349_clk_i memory\[17\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11514_ _05699_ _05714_ _05729_ _05730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_0_81_745 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_81_767 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15282_ _00241_ clknet_leaf_39_clk_i memory\[47\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12494_ _06695_ _06696_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__inv_1
Xclkbuf_leaf_296_clk_i clknet_5_15__leaf_clk_i clknet_leaf_296_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_135_184 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11036__I0 _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14233_ _01272_ clknet_leaf_109_clk_i memory\[12\]\[29\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11445_ _03119_ _05661_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_8
XANTENNA__10815__S _05312_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13281__S0 _02205_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11736__A1 _05676_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07396__S _03437_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14164_ _01203_ clknet_leaf_136_clk_i memory\[7\]\[24\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11376_ _05620_ _00702_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_132_891 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_150_198 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_42_1118 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13115_ _02375_ _02510_ _02511_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_EDGE_ROW_156_Right_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_10327_ _05060_ memory\[46\]\[26\] _05048_ _05061_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14095_ _01134_ clknet_leaf_248_clk_i memory\[63\]\[19\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_13046_ _02358_ _02435_ _02442_ _02443_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__09401__I0 _04189_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10258_ _03137_ _05014_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XTAP_TAPCELL_ROW_167_3592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__07168__A1 net5 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__10550__S _05181_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_128_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10189_ _04975_ _00160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_128_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_234_clk_i clknet_5_15__leaf_clk_i clknet_leaf_234_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__13146__B _02195_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13336__S1 _05779_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_191_1122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_156_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__12839__I1 net49 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_834 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14997_ _02036_ clknet_leaf_64_clk_i memory\[38\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_88_311 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_152_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13948_ _00987_ clknet_leaf_345_clk_i memory\[49\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_117_1237 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_156_1297 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__07715__I0 _03160_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13661__A1 _05654_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12464__A2 _06666_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_89_889 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_92_1285 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_249_clk_i clknet_5_25__leaf_clk_i clknet_leaf_249_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_5_1001 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_53_1258 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13879_ _00918_ clknet_leaf_18_clk_i memory\[39\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11381__S _05616_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_29_422 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_9_1192 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15618_ _00577_ clknet_leaf_322_clk_i memory\[58\]\[6\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_159_799 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__08754__I _03128_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_118_107 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_174_747 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_1067 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12276__I _05791_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_15549_ _00508_ clknet_leaf_333_clk_i memory\[56\]\[1\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08140__I0 _03754_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_84_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_127_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11975__A1 _05753_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09786__S _04751_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_126_151 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09070_ _04366_ _01730_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_167_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_4_522 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08021_ _03787_ memory\[12\]\[17\] _03773_ _03788_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_25_661 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_21_72 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_53_970 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_953 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_112_96 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_71_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_188_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_24_171 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_102_519 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_142_699 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_24_193 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_97_54 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_TAPCELL_ROW_90_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_12_366 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_90_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_97_76 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_187_3968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_187_3979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_EDGE_ROW_123_Right_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_0_750 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_09972_ net72 _04787_ _04860_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_0_772 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_08923_ _04187_ memory\[27\]\[2\] _04286_ _04289_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__12152__A1 _06146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_97_1141 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__10460__S _05131_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_23_1095 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08854_ _04252_ _01628_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07954__I0 _03212_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_34_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_EDGE_ROW_179_Left_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__09026__S _04333_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07805_ _03663_ _01168_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_08785_ _03159_ _04206_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_4
XFILLER_0_19_1109 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_88_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_88_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07736_ _03191_ memory\[63\]\[21\] _03625_ _03627_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_0_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_0_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08865__S _04250_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13652__A1 _05777_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_135_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__07706__I0 _03147_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_49_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_49_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07667_ _03590_ _01103_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_138_928 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09406_ _04544_ _01888_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_164_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_153_92 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_149_276 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09459__I0 _04247_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07598_ _03553_ _01071_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_48_775 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09337_ _04193_ memory\[33\]\[5\] _04502_ _04508_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XPHY_EDGE_ROW_188_Left_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_0_36_959 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_62_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_106_803 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_118_663 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_168_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_129_1119 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09268_ _04471_ _01823_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_62_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_63_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_08219_ _03900_ _01345_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11018__I0 _05064_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12914__I _05683_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09199_ _04191_ memory\[31\]\[4\] _04430_ _04435_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__10635__S _05218_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_69_1298 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_160_452 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11718__A1 _05783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13011__S _02193_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11230_ _03490_ _03750_ _05542_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XANTENNA__08105__S _03830_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09631__I0 _04573_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11161_ _05505_ _00602_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10434__I _05108_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12850__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07944__S _03733_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10112_ _04577_ memory\[44\]\[1\] _04933_ _04935_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_8_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11092_ _05070_ memory\[57\]\[31\] _05434_ _05469_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__13566__S1 _03748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_8_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08198__I0 _03812_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10043_ _04898_ _00091_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14920_ _01959_ clknet_leaf_36_clk_i memory\[36\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_TAPCELL_ROW_145_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_145_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1214 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_11_clk_i_I clknet_5_5__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14851_ _01890_ clknet_leaf_428_clk_i memory\[34\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_98_620 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_106_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_106_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13802_ _00841_ clknet_leaf_207_clk_i memory\[16\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_187_316 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_193_4106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14782_ _01821_ clknet_leaf_426_clk_i memory\[32\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__13643__A1 _05752_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11994_ memory\[16\]\[6\] memory\[17\]\[6\] memory\[18\]\[6\] memory\[19\]\[6\] _05795_
+ _05796_ _06204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_98_664 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_187_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_123_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_13733_ _03098_ _00783_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_303 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__12297__S _06421_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_10945_ _05391_ _00500_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_156_714 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_500 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13664_ memory\[46\]\[31\] memory\[47\]\[31\] _02487_ _03051_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_116_1292 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10876_ _05354_ _00468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_13_1220 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_2_1218 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_15403_ _00362_ clknet_leaf_238_clk_i memory\[51\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__11257__I0 _03334_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12615_ _06480_ _06815_ _06482_ _06816_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__12096__I _05664_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_94_881 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_155_246 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_137_950 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_236_clk_i_I clknet_5_26__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08122__I0 _03806_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13595_ _05660_ _02982_ _05708_ _02983_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_143_408 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_170_205 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_5_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_87_1332 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_171_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_26_447 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15334_ _00293_ clknet_leaf_237_clk_i memory\[4\]\[10\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12546_ _06603_ _06743_ _06745_ _06747_ _06748_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XANTENNA__08673__I1 _03367_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_170_238 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_123_121 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_15265_ _00224_ clknet_leaf_417_clk_i memory\[47\]\[5\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_12477_ _06480_ _06679_ _06482_ _06680_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__12057__S1 _05796_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_152_986 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_169_3621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_14216_ _01255_ clknet_leaf_217_clk_i memory\[12\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__08015__S _03773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_11428_ _05647_ _00727_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_169_3632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15196_ _00155_ clknet_leaf_423_clk_i memory\[45\]\[0\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_50_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12382__A1 _06428_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_349 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_46_1073 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_14147_ _01186_ clknet_leaf_286_clk_i memory\[7\]\[7\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11359_ memory\[61\]\[28\] _03211_ _05602_ _05611_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_120_850 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_158_37 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__13006__S0 _06709_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14078_ _01117_ clknet_leaf_310_clk_i memory\[63\]\[2\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_173_clk_i clknet_5_28__leaf_clk_i clknet_leaf_173_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_20_1224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_13029_ _02216_ _02425_ _02426_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_TAPCELL_ROW_182_3876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__08749__I _03110_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_177_2 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_158_1359 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_83_34 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_08570_ _04086_ _01510_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__08685__S _04146_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__09689__I0 _04633_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_188_clk_i clknet_5_29__leaf_clk_i clknet_leaf_188_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_07521_ memory\[59\]\[17\] _03344_ _03504_ _03512_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_57_1180 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_159_530 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_88_163 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_193_308 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_07452_ _03474_ _01004_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_92_807 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_130_1223 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_230 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_76_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_29_241 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_393 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_111_clk_i clknet_5_23__leaf_clk_i clknet_leaf_111_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_147_758 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_9_647 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_135_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__11248__I0 _03325_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_07383_ _03184_ memory\[8\]\[19\] _03426_ _03436_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_TAPCELL_ROW_44_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_44_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_162_728 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_09122_ _04393_ _04394_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_0_146_279 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_162_739 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09861__I0 _04598_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09053_ _03528_ net72 _04357_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__nand2_4
XFILLER_0_114_132 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_143_975 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_126_clk_i clknet_5_29__leaf_clk_i clknet_leaf_126_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_08004_ _03776_ _01254_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_130_603 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_1152 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_114_154 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_143_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_163_1054 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__13165__A3 _02559_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_41_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__09613__I0 _04625_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__12373__A1 _06155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_13_686 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_438_clk_i_I clknet_5_0__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_861 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__07764__S _03639_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__13548__S1 _02502_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09955_ _04851_ _00050_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_0_580 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__11286__S _05565_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_0_591 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_5_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_08906_ _04279_ _01653_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__10190__S _04969_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_09886_ _04623_ memory\[40\]\[23\] _04811_ _04815_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__07927__I0 _03172_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08837_ _03211_ _04241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA_clkbuf_leaf_185_clk_i_I clknet_5_29__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07552__A1 _03112_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08768_ _04194_ _01600_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_68_804 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_140_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_140_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_07719_ _03166_ memory\[63\]\[13\] _03614_ _03618_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_36_1242 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_95_623 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__11813__I _05677_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__08352__I0 _03762_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_08699_ _03768_ memory\[24\]\[8\] _04146_ _04155_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_135_1189 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_64_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_67_336 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_64_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_137_202 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_32_1117 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_133 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_101_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_10730_ _05277_ _00399_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_TAPCELL_ROW_101_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_83_818 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_36_701 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_94_166 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_870 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_81_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_81_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_94_177 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_10661_ memory\[51\]\[20\] _03186_ _05240_ _05241_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_153_706 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_24_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_24_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_48_594 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_119_972 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12400_ _05655_ _06604_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_13380_ memory\[52\]\[27\] memory\[53\]\[27\] _05716_ _02771_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_63_553 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_10592_ _05047_ memory\[50\]\[20\] _05203_ _05204_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__09852__I0 _04589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_36_778 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__12600__A2 _06800_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_134_942 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1_1262 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_12331_ _06318_ _06531_ _06533_ _06535_ _06536_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_0_35_288 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_12262_ memory\[28\]\[10\] memory\[29\]\[10\] _05915_ _06468_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_50_247 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15050_ _00009_ clknet_leaf_32_clk_i memory\[40\]\[14\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_47_1360 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12364__A1 _06149_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14001_ _01040_ clknet_leaf_165_clk_i memory\[59\]\[21\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_11213_ _05533_ _00626_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__11411__I0 _03350_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_12193_ _05914_ _06395_ _06397_ _06399_ _06400_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
Xclkbuf_leaf_90_clk_i clknet_5_20__leaf_clk_i clknet_leaf_90_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_147_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_TAPCELL_ROW_147_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_31_494 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput41 net41 data_o[10] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__buf_3
XANTENNA__07674__S _03589_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput52 net52 data_o[20] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
X_11144_ _03357_ memory\[58\]\[23\] _05493_ _05497_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
Xoutput63 net63 data_o[30] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_4
XANTENNA__12116__A1 _06322_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_164_3540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_11075_ _05460_ _00561_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_179_1083 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_179_1094 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_125_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_76_1011 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10026_ _04627_ memory\[42\]\[25\] _04883_ _04889_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_14903_ _01942_ clknet_leaf_73_clk_i memory\[35\]\[27\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_76_1033 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_TAPCELL_ROW_160_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__11924__S _05656_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_14834_ _01873_ clknet_leaf_75_clk_i memory\[33\]\[22\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__12419__A2 _06586_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_TAPCELL_ROW_121_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_37_1039 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_76_1099 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_612 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_14765_ _01804_ clknet_leaf_128_clk_i memory\[31\]\[17\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_58_314 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_100 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_11977_ memory\[40\]\[6\] memory\[41\]\[6\] memory\[42\]\[6\] memory\[43\]\[6\] _06186_
+ _05762_ _06187_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_2
XFILLER_0_58_325 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_175_319 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_85_122 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13716_ _03089_ _00775_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_85_144 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_86_667 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_10928_ _05382_ _00492_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_14696_ _01735_ clknet_leaf_168_clk_i memory\[2\]\[12\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_15_1348 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_58_369 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_128_224 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_39_572 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_117_909 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_387_clk_i_I clknet_5_6__leaf_clk_i vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_13647_ memory\[12\]\[31\] memory\[13\]\[31\] _05769_ _03034_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_0_67_892 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_183_352 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_10859_ _05345_ _00460_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__07849__S _03686_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_26_233 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_171_525 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_43_clk_i clknet_5_18__leaf_clk_i clknet_leaf_43_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__08646__I1 _03340_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_147_1016 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_13578_ _02965_ _02966_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_0_48_1102 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_186_1087 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15317_ _00276_ clknet_leaf_263_clk_i memory\[48\]\[25\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_42_737 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_12529_ memory\[32\]\[14\] memory\[33\]\[14\] memory\[34\]\[14\] memory\[35\]\[14\]
+ _06314_ _06454_ _06731_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_0_26_299 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_2_801 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_136_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_125_997 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_48_1157 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_151_260 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_23_962 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_15248_ _00207_ clknet_leaf_154_clk_i memory\[46\]\[20\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_0_151_282 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_140_967 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__13586__S _05773_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_112_658 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__12355__A1 _06276_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__11402__I0 _03342_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_111_135 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_TAPCELL_ROW_184_3905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_58_clk_i clknet_5_17__leaf_clk_i clknet_leaf_58_clk_i vdd vdd vss vss
+ gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_TAPCELL_ROW_184_3916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_15179_ _00138_ clknet_leaf_38_clk_i memory\[44\]\[15\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__09071__I1 memory\[2\]\[8\] vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07584__S _03541_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__07082__I0 _03203_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_123_1060 vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_06952_ _03169_ memory\[14\]\[14\] _03157_ _03170_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_09740_ _04713_ _04736_ vdd vdd vss vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
.ends

