magic
tech gf180mcuD
magscale 1 10
timestamp 1701783334
<< metal1 >>
rect 16818 16718 16830 16770
rect 16882 16767 16894 16770
rect 17378 16767 17390 16770
rect 16882 16721 17390 16767
rect 16882 16718 16894 16721
rect 17378 16718 17390 16721
rect 17442 16718 17454 16770
rect 18162 16718 18174 16770
rect 18226 16767 18238 16770
rect 18834 16767 18846 16770
rect 18226 16721 18846 16767
rect 18226 16718 18238 16721
rect 18834 16718 18846 16721
rect 18898 16718 18910 16770
rect 1344 16490 18592 16524
rect 1344 16438 3370 16490
rect 3422 16438 3474 16490
rect 3526 16438 3578 16490
rect 3630 16438 7682 16490
rect 7734 16438 7786 16490
rect 7838 16438 7890 16490
rect 7942 16438 11994 16490
rect 12046 16438 12098 16490
rect 12150 16438 12202 16490
rect 12254 16438 16306 16490
rect 16358 16438 16410 16490
rect 16462 16438 16514 16490
rect 16566 16438 18592 16490
rect 1344 16404 18592 16438
rect 5966 16322 6018 16334
rect 5966 16258 6018 16270
rect 2706 16158 2718 16210
rect 2770 16158 2782 16210
rect 4050 16158 4062 16210
rect 4114 16158 4126 16210
rect 7646 16098 7698 16110
rect 3154 16046 3166 16098
rect 3218 16046 3230 16098
rect 4946 16046 4958 16098
rect 5010 16046 5022 16098
rect 6626 16046 6638 16098
rect 6690 16046 6702 16098
rect 7646 16034 7698 16046
rect 11006 16098 11058 16110
rect 11006 16034 11058 16046
rect 7086 15986 7138 15998
rect 7086 15922 7138 15934
rect 8766 15986 8818 15998
rect 8766 15922 8818 15934
rect 9662 15986 9714 15998
rect 9662 15922 9714 15934
rect 10334 15986 10386 15998
rect 10334 15922 10386 15934
rect 11678 15986 11730 15998
rect 11678 15922 11730 15934
rect 12350 15986 12402 15998
rect 12350 15922 12402 15934
rect 13134 15986 13186 15998
rect 13134 15922 13186 15934
rect 13694 15986 13746 15998
rect 13694 15922 13746 15934
rect 14366 15986 14418 15998
rect 14366 15922 14418 15934
rect 15038 15986 15090 15998
rect 15038 15922 15090 15934
rect 15710 15986 15762 15998
rect 15710 15922 15762 15934
rect 16942 15986 16994 15998
rect 16942 15922 16994 15934
rect 17390 15986 17442 15998
rect 17390 15922 17442 15934
rect 17838 15986 17890 15998
rect 17838 15922 17890 15934
rect 1710 15874 1762 15886
rect 1710 15810 1762 15822
rect 7982 15874 8034 15886
rect 7982 15810 8034 15822
rect 11342 15874 11394 15886
rect 11342 15810 11394 15822
rect 16382 15874 16434 15886
rect 16382 15810 16434 15822
rect 1344 15706 18752 15740
rect 1344 15654 5526 15706
rect 5578 15654 5630 15706
rect 5682 15654 5734 15706
rect 5786 15654 9838 15706
rect 9890 15654 9942 15706
rect 9994 15654 10046 15706
rect 10098 15654 14150 15706
rect 14202 15654 14254 15706
rect 14306 15654 14358 15706
rect 14410 15654 18462 15706
rect 18514 15654 18566 15706
rect 18618 15654 18670 15706
rect 18722 15654 18752 15706
rect 1344 15620 18752 15654
rect 3614 15538 3666 15550
rect 3614 15474 3666 15486
rect 5630 15538 5682 15550
rect 5630 15474 5682 15486
rect 6302 15538 6354 15550
rect 6302 15474 6354 15486
rect 7422 15538 7474 15550
rect 7422 15474 7474 15486
rect 8318 15538 8370 15550
rect 8318 15474 8370 15486
rect 10782 15538 10834 15550
rect 10782 15474 10834 15486
rect 17726 15538 17778 15550
rect 17726 15474 17778 15486
rect 18174 15538 18226 15550
rect 18174 15474 18226 15486
rect 1710 15426 1762 15438
rect 1710 15362 1762 15374
rect 1344 14922 18592 14956
rect 1344 14870 3370 14922
rect 3422 14870 3474 14922
rect 3526 14870 3578 14922
rect 3630 14870 7682 14922
rect 7734 14870 7786 14922
rect 7838 14870 7890 14922
rect 7942 14870 11994 14922
rect 12046 14870 12098 14922
rect 12150 14870 12202 14922
rect 12254 14870 16306 14922
rect 16358 14870 16410 14922
rect 16462 14870 16514 14922
rect 16566 14870 18592 14922
rect 1344 14836 18592 14870
rect 10434 14478 10446 14530
rect 10498 14478 10510 14530
rect 6178 14366 6190 14418
rect 6242 14366 6254 14418
rect 1710 14306 1762 14318
rect 1710 14242 1762 14254
rect 1344 14138 18752 14172
rect 1344 14086 5526 14138
rect 5578 14086 5630 14138
rect 5682 14086 5734 14138
rect 5786 14086 9838 14138
rect 9890 14086 9942 14138
rect 9994 14086 10046 14138
rect 10098 14086 14150 14138
rect 14202 14086 14254 14138
rect 14306 14086 14358 14138
rect 14410 14086 18462 14138
rect 18514 14086 18566 14138
rect 18618 14086 18670 14138
rect 18722 14086 18752 14138
rect 1344 14052 18752 14086
rect 1710 13858 1762 13870
rect 1710 13794 1762 13806
rect 1344 13354 18592 13388
rect 1344 13302 3370 13354
rect 3422 13302 3474 13354
rect 3526 13302 3578 13354
rect 3630 13302 7682 13354
rect 7734 13302 7786 13354
rect 7838 13302 7890 13354
rect 7942 13302 11994 13354
rect 12046 13302 12098 13354
rect 12150 13302 12202 13354
rect 12254 13302 16306 13354
rect 16358 13302 16410 13354
rect 16462 13302 16514 13354
rect 16566 13302 18592 13354
rect 1344 13268 18592 13302
rect 1344 12570 18752 12604
rect 1344 12518 5526 12570
rect 5578 12518 5630 12570
rect 5682 12518 5734 12570
rect 5786 12518 9838 12570
rect 9890 12518 9942 12570
rect 9994 12518 10046 12570
rect 10098 12518 14150 12570
rect 14202 12518 14254 12570
rect 14306 12518 14358 12570
rect 14410 12518 18462 12570
rect 18514 12518 18566 12570
rect 18618 12518 18670 12570
rect 18722 12518 18752 12570
rect 1344 12484 18752 12518
rect 1710 12290 1762 12302
rect 1710 12226 1762 12238
rect 9886 12290 9938 12302
rect 9886 12226 9938 12238
rect 10334 12290 10386 12302
rect 10334 12226 10386 12238
rect 6178 12126 6190 12178
rect 6242 12126 6254 12178
rect 6850 12014 6862 12066
rect 6914 12014 6926 12066
rect 8978 12014 8990 12066
rect 9042 12014 9054 12066
rect 5742 11954 5794 11966
rect 5742 11890 5794 11902
rect 9774 11954 9826 11966
rect 9774 11890 9826 11902
rect 10222 11954 10274 11966
rect 10222 11890 10274 11902
rect 1344 11786 18592 11820
rect 1344 11734 3370 11786
rect 3422 11734 3474 11786
rect 3526 11734 3578 11786
rect 3630 11734 7682 11786
rect 7734 11734 7786 11786
rect 7838 11734 7890 11786
rect 7942 11734 11994 11786
rect 12046 11734 12098 11786
rect 12150 11734 12202 11786
rect 12254 11734 16306 11786
rect 16358 11734 16410 11786
rect 16462 11734 16514 11786
rect 16566 11734 18592 11786
rect 1344 11700 18592 11734
rect 5182 11394 5234 11406
rect 1810 11342 1822 11394
rect 1874 11342 1886 11394
rect 6402 11342 6414 11394
rect 6466 11342 6478 11394
rect 5182 11330 5234 11342
rect 5742 11282 5794 11294
rect 5742 11218 5794 11230
rect 6078 11282 6130 11294
rect 10434 11230 10446 11282
rect 10498 11230 10510 11282
rect 6078 11218 6130 11230
rect 2046 11170 2098 11182
rect 2046 11106 2098 11118
rect 2494 11170 2546 11182
rect 2494 11106 2546 11118
rect 1344 11002 18752 11036
rect 1344 10950 5526 11002
rect 5578 10950 5630 11002
rect 5682 10950 5734 11002
rect 5786 10950 9838 11002
rect 9890 10950 9942 11002
rect 9994 10950 10046 11002
rect 10098 10950 14150 11002
rect 14202 10950 14254 11002
rect 14306 10950 14358 11002
rect 14410 10950 18462 11002
rect 18514 10950 18566 11002
rect 18618 10950 18670 11002
rect 18722 10950 18752 11002
rect 1344 10916 18752 10950
rect 9102 10834 9154 10846
rect 8306 10782 8318 10834
rect 8370 10782 8382 10834
rect 9102 10770 9154 10782
rect 1710 10722 1762 10734
rect 1710 10658 1762 10670
rect 9998 10722 10050 10734
rect 12574 10722 12626 10734
rect 11778 10670 11790 10722
rect 11842 10670 11854 10722
rect 9998 10658 10050 10670
rect 12574 10658 12626 10670
rect 5406 10610 5458 10622
rect 9886 10610 9938 10622
rect 12462 10610 12514 10622
rect 5954 10558 5966 10610
rect 6018 10558 6030 10610
rect 11666 10558 11678 10610
rect 11730 10558 11742 10610
rect 5406 10546 5458 10558
rect 9886 10546 9938 10558
rect 12462 10546 12514 10558
rect 10894 10498 10946 10510
rect 10894 10434 10946 10446
rect 9998 10386 10050 10398
rect 9998 10322 10050 10334
rect 11230 10386 11282 10398
rect 11230 10322 11282 10334
rect 12574 10386 12626 10398
rect 12574 10322 12626 10334
rect 1344 10218 18592 10252
rect 1344 10166 3370 10218
rect 3422 10166 3474 10218
rect 3526 10166 3578 10218
rect 3630 10166 7682 10218
rect 7734 10166 7786 10218
rect 7838 10166 7890 10218
rect 7942 10166 11994 10218
rect 12046 10166 12098 10218
rect 12150 10166 12202 10218
rect 12254 10166 16306 10218
rect 16358 10166 16410 10218
rect 16462 10166 16514 10218
rect 16566 10166 18592 10218
rect 1344 10132 18592 10166
rect 12238 10050 12290 10062
rect 12238 9986 12290 9998
rect 12450 9886 12462 9938
rect 12514 9886 12526 9938
rect 13358 9826 13410 9838
rect 7634 9774 7646 9826
rect 7698 9774 7710 9826
rect 8082 9774 8094 9826
rect 8146 9774 8158 9826
rect 11890 9774 11902 9826
rect 11954 9774 11966 9826
rect 13358 9762 13410 9774
rect 10670 9714 10722 9726
rect 8194 9662 8206 9714
rect 8258 9662 8270 9714
rect 10670 9650 10722 9662
rect 12462 9714 12514 9726
rect 12462 9650 12514 9662
rect 13582 9714 13634 9726
rect 13582 9650 13634 9662
rect 13694 9714 13746 9726
rect 13694 9650 13746 9662
rect 7422 9602 7474 9614
rect 7422 9538 7474 9550
rect 11118 9602 11170 9614
rect 11118 9538 11170 9550
rect 1344 9434 18752 9468
rect 1344 9382 5526 9434
rect 5578 9382 5630 9434
rect 5682 9382 5734 9434
rect 5786 9382 9838 9434
rect 9890 9382 9942 9434
rect 9994 9382 10046 9434
rect 10098 9382 14150 9434
rect 14202 9382 14254 9434
rect 14306 9382 14358 9434
rect 14410 9382 18462 9434
rect 18514 9382 18566 9434
rect 18618 9382 18670 9434
rect 18722 9382 18752 9434
rect 1344 9348 18752 9382
rect 9102 9266 9154 9278
rect 8306 9214 8318 9266
rect 8370 9214 8382 9266
rect 9102 9202 9154 9214
rect 9662 9266 9714 9278
rect 11778 9214 11790 9266
rect 11842 9214 11854 9266
rect 9662 9202 9714 9214
rect 17838 9154 17890 9166
rect 10322 9102 10334 9154
rect 10386 9102 10398 9154
rect 10546 9102 10558 9154
rect 10610 9102 10622 9154
rect 11330 9102 11342 9154
rect 11394 9102 11406 9154
rect 12786 9102 12798 9154
rect 12850 9102 12862 9154
rect 13458 9102 13470 9154
rect 13522 9102 13534 9154
rect 17838 9090 17890 9102
rect 5630 9042 5682 9054
rect 9998 9042 10050 9054
rect 12350 9042 12402 9054
rect 18174 9042 18226 9054
rect 6066 8990 6078 9042
rect 6130 8990 6142 9042
rect 11778 8990 11790 9042
rect 11842 8990 11854 9042
rect 13346 8990 13358 9042
rect 13410 8990 13422 9042
rect 13906 8990 13918 9042
rect 13970 8990 13982 9042
rect 14690 8990 14702 9042
rect 14754 8990 14766 9042
rect 5630 8978 5682 8990
rect 9998 8978 10050 8990
rect 12350 8978 12402 8990
rect 18174 8978 18226 8990
rect 17614 8930 17666 8942
rect 17614 8866 17666 8878
rect 14478 8818 14530 8830
rect 14478 8754 14530 8766
rect 1344 8650 18592 8684
rect 1344 8598 3370 8650
rect 3422 8598 3474 8650
rect 3526 8598 3578 8650
rect 3630 8598 7682 8650
rect 7734 8598 7786 8650
rect 7838 8598 7890 8650
rect 7942 8598 11994 8650
rect 12046 8598 12098 8650
rect 12150 8598 12202 8650
rect 12254 8598 16306 8650
rect 16358 8598 16410 8650
rect 16462 8598 16514 8650
rect 16566 8598 18592 8650
rect 1344 8564 18592 8598
rect 6626 8318 6638 8370
rect 6690 8318 6702 8370
rect 12674 8318 12686 8370
rect 12738 8318 12750 8370
rect 10434 8206 10446 8258
rect 10498 8206 10510 8258
rect 12562 8206 12574 8258
rect 12626 8206 12638 8258
rect 1710 8146 1762 8158
rect 1710 8082 1762 8094
rect 12910 8146 12962 8158
rect 12910 8082 12962 8094
rect 17166 8146 17218 8158
rect 17166 8082 17218 8094
rect 17502 8146 17554 8158
rect 17502 8082 17554 8094
rect 17838 8146 17890 8158
rect 17838 8082 17890 8094
rect 18174 8146 18226 8158
rect 18174 8082 18226 8094
rect 2046 8034 2098 8046
rect 2046 7970 2098 7982
rect 2382 8034 2434 8046
rect 2382 7970 2434 7982
rect 1344 7866 18752 7900
rect 1344 7814 5526 7866
rect 5578 7814 5630 7866
rect 5682 7814 5734 7866
rect 5786 7814 9838 7866
rect 9890 7814 9942 7866
rect 9994 7814 10046 7866
rect 10098 7814 14150 7866
rect 14202 7814 14254 7866
rect 14306 7814 14358 7866
rect 14410 7814 18462 7866
rect 18514 7814 18566 7866
rect 18618 7814 18670 7866
rect 18722 7814 18752 7866
rect 1344 7780 18752 7814
rect 1822 7698 1874 7710
rect 1822 7634 1874 7646
rect 13806 7698 13858 7710
rect 13806 7634 13858 7646
rect 18286 7698 18338 7710
rect 18286 7634 18338 7646
rect 11118 7586 11170 7598
rect 7410 7534 7422 7586
rect 7474 7534 7486 7586
rect 8978 7534 8990 7586
rect 9042 7534 9054 7586
rect 11118 7522 11170 7534
rect 13134 7586 13186 7598
rect 13134 7522 13186 7534
rect 8430 7474 8482 7486
rect 17726 7474 17778 7486
rect 7298 7422 7310 7474
rect 7362 7422 7374 7474
rect 9874 7422 9886 7474
rect 9938 7422 9950 7474
rect 10546 7422 10558 7474
rect 10610 7422 10622 7474
rect 14354 7422 14366 7474
rect 14418 7422 14430 7474
rect 8430 7410 8482 7422
rect 17726 7410 17778 7422
rect 8306 7310 8318 7362
rect 8370 7310 8382 7362
rect 9986 7310 9998 7362
rect 10050 7310 10062 7362
rect 10222 7250 10274 7262
rect 10222 7186 10274 7198
rect 1344 7082 18592 7116
rect 1344 7030 3370 7082
rect 3422 7030 3474 7082
rect 3526 7030 3578 7082
rect 3630 7030 7682 7082
rect 7734 7030 7786 7082
rect 7838 7030 7890 7082
rect 7942 7030 11994 7082
rect 12046 7030 12098 7082
rect 12150 7030 12202 7082
rect 12254 7030 16306 7082
rect 16358 7030 16410 7082
rect 16462 7030 16514 7082
rect 16566 7030 18592 7082
rect 1344 6996 18592 7030
rect 12574 6690 12626 6702
rect 8194 6638 8206 6690
rect 8258 6638 8270 6690
rect 10210 6638 10222 6690
rect 10274 6638 10286 6690
rect 12574 6626 12626 6638
rect 12910 6690 12962 6702
rect 12910 6626 12962 6638
rect 8766 6578 8818 6590
rect 8766 6514 8818 6526
rect 10782 6578 10834 6590
rect 10782 6514 10834 6526
rect 12686 6578 12738 6590
rect 12686 6514 12738 6526
rect 1822 6466 1874 6478
rect 9650 6414 9662 6466
rect 9714 6414 9726 6466
rect 1822 6402 1874 6414
rect 1344 6298 18752 6332
rect 1344 6246 5526 6298
rect 5578 6246 5630 6298
rect 5682 6246 5734 6298
rect 5786 6246 9838 6298
rect 9890 6246 9942 6298
rect 9994 6246 10046 6298
rect 10098 6246 14150 6298
rect 14202 6246 14254 6298
rect 14306 6246 14358 6298
rect 14410 6246 18462 6298
rect 18514 6246 18566 6298
rect 18618 6246 18670 6298
rect 18722 6246 18752 6298
rect 1344 6212 18752 6246
rect 10334 6130 10386 6142
rect 13570 6078 13582 6130
rect 13634 6078 13646 6130
rect 10334 6066 10386 6078
rect 1710 6018 1762 6030
rect 10222 6018 10274 6030
rect 7074 5966 7086 6018
rect 7138 5966 7150 6018
rect 8754 5966 8766 6018
rect 8818 5966 8830 6018
rect 1710 5954 1762 5966
rect 10222 5954 10274 5966
rect 12014 6018 12066 6030
rect 14466 5966 14478 6018
rect 14530 5966 14542 6018
rect 12014 5954 12066 5966
rect 7746 5854 7758 5906
rect 7810 5854 7822 5906
rect 8082 5854 8094 5906
rect 8146 5854 8158 5906
rect 12562 5854 12574 5906
rect 12626 5854 12638 5906
rect 14578 5854 14590 5906
rect 14642 5854 14654 5906
rect 2270 5794 2322 5806
rect 2270 5730 2322 5742
rect 2718 5794 2770 5806
rect 17614 5794 17666 5806
rect 8306 5742 8318 5794
rect 8370 5742 8382 5794
rect 2718 5730 2770 5742
rect 17614 5730 17666 5742
rect 18286 5794 18338 5806
rect 18286 5730 18338 5742
rect 10446 5682 10498 5694
rect 10446 5618 10498 5630
rect 1344 5514 18592 5548
rect 1344 5462 3370 5514
rect 3422 5462 3474 5514
rect 3526 5462 3578 5514
rect 3630 5462 7682 5514
rect 7734 5462 7786 5514
rect 7838 5462 7890 5514
rect 7942 5462 11994 5514
rect 12046 5462 12098 5514
rect 12150 5462 12202 5514
rect 12254 5462 16306 5514
rect 16358 5462 16410 5514
rect 16462 5462 16514 5514
rect 16566 5462 18592 5514
rect 1344 5428 18592 5462
rect 11118 5346 11170 5358
rect 11118 5282 11170 5294
rect 1710 5122 1762 5134
rect 1710 5058 1762 5070
rect 3614 5122 3666 5134
rect 11006 5122 11058 5134
rect 9538 5070 9550 5122
rect 9602 5070 9614 5122
rect 10322 5070 10334 5122
rect 10386 5070 10398 5122
rect 3614 5058 3666 5070
rect 11006 5058 11058 5070
rect 16718 5122 16770 5134
rect 16718 5058 16770 5070
rect 17166 5122 17218 5134
rect 17166 5058 17218 5070
rect 18174 5122 18226 5134
rect 18174 5058 18226 5070
rect 2046 5010 2098 5022
rect 17838 5010 17890 5022
rect 9650 4958 9662 5010
rect 9714 4958 9726 5010
rect 2046 4946 2098 4958
rect 17838 4946 17890 4958
rect 2382 4898 2434 4910
rect 2382 4834 2434 4846
rect 3166 4898 3218 4910
rect 3166 4834 3218 4846
rect 15598 4898 15650 4910
rect 15598 4834 15650 4846
rect 17614 4898 17666 4910
rect 17614 4834 17666 4846
rect 1344 4730 18752 4764
rect 1344 4678 5526 4730
rect 5578 4678 5630 4730
rect 5682 4678 5734 4730
rect 5786 4678 9838 4730
rect 9890 4678 9942 4730
rect 9994 4678 10046 4730
rect 10098 4678 14150 4730
rect 14202 4678 14254 4730
rect 14306 4678 14358 4730
rect 14410 4678 18462 4730
rect 18514 4678 18566 4730
rect 18618 4678 18670 4730
rect 18722 4678 18752 4730
rect 1344 4644 18752 4678
rect 2046 4562 2098 4574
rect 2046 4498 2098 4510
rect 2718 4562 2770 4574
rect 2718 4498 2770 4510
rect 5966 4562 6018 4574
rect 5966 4498 6018 4510
rect 15710 4562 15762 4574
rect 15710 4498 15762 4510
rect 16494 4562 16546 4574
rect 16494 4498 16546 4510
rect 3054 4450 3106 4462
rect 3054 4386 3106 4398
rect 17726 4450 17778 4462
rect 17726 4386 17778 4398
rect 1710 4338 1762 4350
rect 1710 4274 1762 4286
rect 2382 4338 2434 4350
rect 2382 4274 2434 4286
rect 5630 4338 5682 4350
rect 16830 4338 16882 4350
rect 15922 4286 15934 4338
rect 15986 4286 15998 4338
rect 17938 4286 17950 4338
rect 18002 4286 18014 4338
rect 5630 4274 5682 4286
rect 16830 4274 16882 4286
rect 3838 4226 3890 4238
rect 3838 4162 3890 4174
rect 4398 4226 4450 4238
rect 4398 4162 4450 4174
rect 4846 4226 4898 4238
rect 4846 4162 4898 4174
rect 5406 4226 5458 4238
rect 5406 4162 5458 4174
rect 6414 4226 6466 4238
rect 6414 4162 6466 4174
rect 6974 4226 7026 4238
rect 6974 4162 7026 4174
rect 7646 4226 7698 4238
rect 7646 4162 7698 4174
rect 8094 4226 8146 4238
rect 8094 4162 8146 4174
rect 8654 4226 8706 4238
rect 8654 4162 8706 4174
rect 9102 4226 9154 4238
rect 9102 4162 9154 4174
rect 10110 4226 10162 4238
rect 10110 4162 10162 4174
rect 10782 4226 10834 4238
rect 10782 4162 10834 4174
rect 11454 4226 11506 4238
rect 11454 4162 11506 4174
rect 13582 4226 13634 4238
rect 13582 4162 13634 4174
rect 14254 4226 14306 4238
rect 14254 4162 14306 4174
rect 14926 4226 14978 4238
rect 14926 4162 14978 4174
rect 15486 4226 15538 4238
rect 15486 4162 15538 4174
rect 1344 3946 18592 3980
rect 1344 3894 3370 3946
rect 3422 3894 3474 3946
rect 3526 3894 3578 3946
rect 3630 3894 7682 3946
rect 7734 3894 7786 3946
rect 7838 3894 7890 3946
rect 7942 3894 11994 3946
rect 12046 3894 12098 3946
rect 12150 3894 12202 3946
rect 12254 3894 16306 3946
rect 16358 3894 16410 3946
rect 16462 3894 16514 3946
rect 16566 3894 18592 3946
rect 1344 3860 18592 3894
rect 1934 3554 1986 3566
rect 11006 3554 11058 3566
rect 12686 3554 12738 3566
rect 15486 3554 15538 3566
rect 2706 3502 2718 3554
rect 2770 3502 2782 3554
rect 3378 3502 3390 3554
rect 3442 3502 3454 3554
rect 4050 3502 4062 3554
rect 4114 3502 4126 3554
rect 4722 3502 4734 3554
rect 4786 3502 4798 3554
rect 5842 3502 5854 3554
rect 5906 3502 5918 3554
rect 6514 3502 6526 3554
rect 6578 3502 6590 3554
rect 7186 3502 7198 3554
rect 7250 3502 7262 3554
rect 7858 3502 7870 3554
rect 7922 3502 7934 3554
rect 8642 3502 8654 3554
rect 8706 3502 8718 3554
rect 9874 3502 9886 3554
rect 9938 3502 9950 3554
rect 10546 3502 10558 3554
rect 10610 3502 10622 3554
rect 11890 3502 11902 3554
rect 11954 3502 11966 3554
rect 13346 3502 13358 3554
rect 13410 3502 13422 3554
rect 14690 3502 14702 3554
rect 14754 3502 14766 3554
rect 16034 3502 16046 3554
rect 16098 3502 16110 3554
rect 17154 3502 17166 3554
rect 17218 3502 17230 3554
rect 1934 3490 1986 3502
rect 11006 3490 11058 3502
rect 12686 3490 12738 3502
rect 15486 3490 15538 3502
rect 2270 3442 2322 3454
rect 2270 3378 2322 3390
rect 4958 3442 5010 3454
rect 4958 3378 5010 3390
rect 8430 3442 8482 3454
rect 8430 3378 8482 3390
rect 9662 3442 9714 3454
rect 9662 3378 9714 3390
rect 11342 3442 11394 3454
rect 11342 3378 11394 3390
rect 11678 3442 11730 3454
rect 11678 3378 11730 3390
rect 13134 3442 13186 3454
rect 13134 3378 13186 3390
rect 14142 3442 14194 3454
rect 14142 3378 14194 3390
rect 14478 3442 14530 3454
rect 14478 3378 14530 3390
rect 15150 3442 15202 3454
rect 15150 3378 15202 3390
rect 15822 3442 15874 3454
rect 15822 3378 15874 3390
rect 16942 3442 16994 3454
rect 16942 3378 16994 3390
rect 17614 3442 17666 3454
rect 17614 3378 17666 3390
rect 17950 3442 18002 3454
rect 17950 3378 18002 3390
rect 2942 3330 2994 3342
rect 2942 3266 2994 3278
rect 3614 3330 3666 3342
rect 6078 3330 6130 3342
rect 4274 3278 4286 3330
rect 4338 3278 4350 3330
rect 3614 3266 3666 3278
rect 6078 3266 6130 3278
rect 6750 3330 6802 3342
rect 6750 3266 6802 3278
rect 7422 3330 7474 3342
rect 7422 3266 7474 3278
rect 8094 3330 8146 3342
rect 8094 3266 8146 3278
rect 10334 3330 10386 3342
rect 10334 3266 10386 3278
rect 13806 3330 13858 3342
rect 13806 3266 13858 3278
rect 1344 3162 18752 3196
rect 1344 3110 5526 3162
rect 5578 3110 5630 3162
rect 5682 3110 5734 3162
rect 5786 3110 9838 3162
rect 9890 3110 9942 3162
rect 9994 3110 10046 3162
rect 10098 3110 14150 3162
rect 14202 3110 14254 3162
rect 14306 3110 14358 3162
rect 14410 3110 18462 3162
rect 18514 3110 18566 3162
rect 18618 3110 18670 3162
rect 18722 3110 18752 3162
rect 1344 3076 18752 3110
rect 16818 2942 16830 2994
rect 16882 2991 16894 2994
rect 17490 2991 17502 2994
rect 16882 2945 17502 2991
rect 16882 2942 16894 2945
rect 17490 2942 17502 2945
rect 17554 2991 17566 2994
rect 17938 2991 17950 2994
rect 17554 2945 17950 2991
rect 17554 2942 17566 2945
rect 17938 2942 17950 2945
rect 18002 2942 18014 2994
<< via1 >>
rect 16830 16718 16882 16770
rect 17390 16718 17442 16770
rect 18174 16718 18226 16770
rect 18846 16718 18898 16770
rect 3370 16438 3422 16490
rect 3474 16438 3526 16490
rect 3578 16438 3630 16490
rect 7682 16438 7734 16490
rect 7786 16438 7838 16490
rect 7890 16438 7942 16490
rect 11994 16438 12046 16490
rect 12098 16438 12150 16490
rect 12202 16438 12254 16490
rect 16306 16438 16358 16490
rect 16410 16438 16462 16490
rect 16514 16438 16566 16490
rect 5966 16270 6018 16322
rect 2718 16158 2770 16210
rect 4062 16158 4114 16210
rect 3166 16046 3218 16098
rect 4958 16046 5010 16098
rect 6638 16046 6690 16098
rect 7646 16046 7698 16098
rect 11006 16046 11058 16098
rect 7086 15934 7138 15986
rect 8766 15934 8818 15986
rect 9662 15934 9714 15986
rect 10334 15934 10386 15986
rect 11678 15934 11730 15986
rect 12350 15934 12402 15986
rect 13134 15934 13186 15986
rect 13694 15934 13746 15986
rect 14366 15934 14418 15986
rect 15038 15934 15090 15986
rect 15710 15934 15762 15986
rect 16942 15934 16994 15986
rect 17390 15934 17442 15986
rect 17838 15934 17890 15986
rect 1710 15822 1762 15874
rect 7982 15822 8034 15874
rect 11342 15822 11394 15874
rect 16382 15822 16434 15874
rect 5526 15654 5578 15706
rect 5630 15654 5682 15706
rect 5734 15654 5786 15706
rect 9838 15654 9890 15706
rect 9942 15654 9994 15706
rect 10046 15654 10098 15706
rect 14150 15654 14202 15706
rect 14254 15654 14306 15706
rect 14358 15654 14410 15706
rect 18462 15654 18514 15706
rect 18566 15654 18618 15706
rect 18670 15654 18722 15706
rect 3614 15486 3666 15538
rect 5630 15486 5682 15538
rect 6302 15486 6354 15538
rect 7422 15486 7474 15538
rect 8318 15486 8370 15538
rect 10782 15486 10834 15538
rect 17726 15486 17778 15538
rect 18174 15486 18226 15538
rect 1710 15374 1762 15426
rect 3370 14870 3422 14922
rect 3474 14870 3526 14922
rect 3578 14870 3630 14922
rect 7682 14870 7734 14922
rect 7786 14870 7838 14922
rect 7890 14870 7942 14922
rect 11994 14870 12046 14922
rect 12098 14870 12150 14922
rect 12202 14870 12254 14922
rect 16306 14870 16358 14922
rect 16410 14870 16462 14922
rect 16514 14870 16566 14922
rect 10446 14478 10498 14530
rect 6190 14366 6242 14418
rect 1710 14254 1762 14306
rect 5526 14086 5578 14138
rect 5630 14086 5682 14138
rect 5734 14086 5786 14138
rect 9838 14086 9890 14138
rect 9942 14086 9994 14138
rect 10046 14086 10098 14138
rect 14150 14086 14202 14138
rect 14254 14086 14306 14138
rect 14358 14086 14410 14138
rect 18462 14086 18514 14138
rect 18566 14086 18618 14138
rect 18670 14086 18722 14138
rect 1710 13806 1762 13858
rect 3370 13302 3422 13354
rect 3474 13302 3526 13354
rect 3578 13302 3630 13354
rect 7682 13302 7734 13354
rect 7786 13302 7838 13354
rect 7890 13302 7942 13354
rect 11994 13302 12046 13354
rect 12098 13302 12150 13354
rect 12202 13302 12254 13354
rect 16306 13302 16358 13354
rect 16410 13302 16462 13354
rect 16514 13302 16566 13354
rect 5526 12518 5578 12570
rect 5630 12518 5682 12570
rect 5734 12518 5786 12570
rect 9838 12518 9890 12570
rect 9942 12518 9994 12570
rect 10046 12518 10098 12570
rect 14150 12518 14202 12570
rect 14254 12518 14306 12570
rect 14358 12518 14410 12570
rect 18462 12518 18514 12570
rect 18566 12518 18618 12570
rect 18670 12518 18722 12570
rect 1710 12238 1762 12290
rect 9886 12238 9938 12290
rect 10334 12238 10386 12290
rect 6190 12126 6242 12178
rect 6862 12014 6914 12066
rect 8990 12014 9042 12066
rect 5742 11902 5794 11954
rect 9774 11902 9826 11954
rect 10222 11902 10274 11954
rect 3370 11734 3422 11786
rect 3474 11734 3526 11786
rect 3578 11734 3630 11786
rect 7682 11734 7734 11786
rect 7786 11734 7838 11786
rect 7890 11734 7942 11786
rect 11994 11734 12046 11786
rect 12098 11734 12150 11786
rect 12202 11734 12254 11786
rect 16306 11734 16358 11786
rect 16410 11734 16462 11786
rect 16514 11734 16566 11786
rect 1822 11342 1874 11394
rect 5182 11342 5234 11394
rect 6414 11342 6466 11394
rect 5742 11230 5794 11282
rect 6078 11230 6130 11282
rect 10446 11230 10498 11282
rect 2046 11118 2098 11170
rect 2494 11118 2546 11170
rect 5526 10950 5578 11002
rect 5630 10950 5682 11002
rect 5734 10950 5786 11002
rect 9838 10950 9890 11002
rect 9942 10950 9994 11002
rect 10046 10950 10098 11002
rect 14150 10950 14202 11002
rect 14254 10950 14306 11002
rect 14358 10950 14410 11002
rect 18462 10950 18514 11002
rect 18566 10950 18618 11002
rect 18670 10950 18722 11002
rect 8318 10782 8370 10834
rect 9102 10782 9154 10834
rect 1710 10670 1762 10722
rect 9998 10670 10050 10722
rect 11790 10670 11842 10722
rect 12574 10670 12626 10722
rect 5406 10558 5458 10610
rect 5966 10558 6018 10610
rect 9886 10558 9938 10610
rect 11678 10558 11730 10610
rect 12462 10558 12514 10610
rect 10894 10446 10946 10498
rect 9998 10334 10050 10386
rect 11230 10334 11282 10386
rect 12574 10334 12626 10386
rect 3370 10166 3422 10218
rect 3474 10166 3526 10218
rect 3578 10166 3630 10218
rect 7682 10166 7734 10218
rect 7786 10166 7838 10218
rect 7890 10166 7942 10218
rect 11994 10166 12046 10218
rect 12098 10166 12150 10218
rect 12202 10166 12254 10218
rect 16306 10166 16358 10218
rect 16410 10166 16462 10218
rect 16514 10166 16566 10218
rect 12238 9998 12290 10050
rect 12462 9886 12514 9938
rect 7646 9774 7698 9826
rect 8094 9774 8146 9826
rect 11902 9774 11954 9826
rect 13358 9774 13410 9826
rect 8206 9662 8258 9714
rect 10670 9662 10722 9714
rect 12462 9662 12514 9714
rect 13582 9662 13634 9714
rect 13694 9662 13746 9714
rect 7422 9550 7474 9602
rect 11118 9550 11170 9602
rect 5526 9382 5578 9434
rect 5630 9382 5682 9434
rect 5734 9382 5786 9434
rect 9838 9382 9890 9434
rect 9942 9382 9994 9434
rect 10046 9382 10098 9434
rect 14150 9382 14202 9434
rect 14254 9382 14306 9434
rect 14358 9382 14410 9434
rect 18462 9382 18514 9434
rect 18566 9382 18618 9434
rect 18670 9382 18722 9434
rect 8318 9214 8370 9266
rect 9102 9214 9154 9266
rect 9662 9214 9714 9266
rect 11790 9214 11842 9266
rect 10334 9102 10386 9154
rect 10558 9102 10610 9154
rect 11342 9102 11394 9154
rect 12798 9102 12850 9154
rect 13470 9102 13522 9154
rect 17838 9102 17890 9154
rect 5630 8990 5682 9042
rect 6078 8990 6130 9042
rect 9998 8990 10050 9042
rect 11790 8990 11842 9042
rect 12350 8990 12402 9042
rect 13358 8990 13410 9042
rect 13918 8990 13970 9042
rect 14702 8990 14754 9042
rect 18174 8990 18226 9042
rect 17614 8878 17666 8930
rect 14478 8766 14530 8818
rect 3370 8598 3422 8650
rect 3474 8598 3526 8650
rect 3578 8598 3630 8650
rect 7682 8598 7734 8650
rect 7786 8598 7838 8650
rect 7890 8598 7942 8650
rect 11994 8598 12046 8650
rect 12098 8598 12150 8650
rect 12202 8598 12254 8650
rect 16306 8598 16358 8650
rect 16410 8598 16462 8650
rect 16514 8598 16566 8650
rect 6638 8318 6690 8370
rect 12686 8318 12738 8370
rect 10446 8206 10498 8258
rect 12574 8206 12626 8258
rect 1710 8094 1762 8146
rect 12910 8094 12962 8146
rect 17166 8094 17218 8146
rect 17502 8094 17554 8146
rect 17838 8094 17890 8146
rect 18174 8094 18226 8146
rect 2046 7982 2098 8034
rect 2382 7982 2434 8034
rect 5526 7814 5578 7866
rect 5630 7814 5682 7866
rect 5734 7814 5786 7866
rect 9838 7814 9890 7866
rect 9942 7814 9994 7866
rect 10046 7814 10098 7866
rect 14150 7814 14202 7866
rect 14254 7814 14306 7866
rect 14358 7814 14410 7866
rect 18462 7814 18514 7866
rect 18566 7814 18618 7866
rect 18670 7814 18722 7866
rect 1822 7646 1874 7698
rect 13806 7646 13858 7698
rect 18286 7646 18338 7698
rect 7422 7534 7474 7586
rect 8990 7534 9042 7586
rect 11118 7534 11170 7586
rect 13134 7534 13186 7586
rect 7310 7422 7362 7474
rect 8430 7422 8482 7474
rect 9886 7422 9938 7474
rect 10558 7422 10610 7474
rect 14366 7422 14418 7474
rect 17726 7422 17778 7474
rect 8318 7310 8370 7362
rect 9998 7310 10050 7362
rect 10222 7198 10274 7250
rect 3370 7030 3422 7082
rect 3474 7030 3526 7082
rect 3578 7030 3630 7082
rect 7682 7030 7734 7082
rect 7786 7030 7838 7082
rect 7890 7030 7942 7082
rect 11994 7030 12046 7082
rect 12098 7030 12150 7082
rect 12202 7030 12254 7082
rect 16306 7030 16358 7082
rect 16410 7030 16462 7082
rect 16514 7030 16566 7082
rect 8206 6638 8258 6690
rect 10222 6638 10274 6690
rect 12574 6638 12626 6690
rect 12910 6638 12962 6690
rect 8766 6526 8818 6578
rect 10782 6526 10834 6578
rect 12686 6526 12738 6578
rect 1822 6414 1874 6466
rect 9662 6414 9714 6466
rect 5526 6246 5578 6298
rect 5630 6246 5682 6298
rect 5734 6246 5786 6298
rect 9838 6246 9890 6298
rect 9942 6246 9994 6298
rect 10046 6246 10098 6298
rect 14150 6246 14202 6298
rect 14254 6246 14306 6298
rect 14358 6246 14410 6298
rect 18462 6246 18514 6298
rect 18566 6246 18618 6298
rect 18670 6246 18722 6298
rect 10334 6078 10386 6130
rect 13582 6078 13634 6130
rect 1710 5966 1762 6018
rect 7086 5966 7138 6018
rect 8766 5966 8818 6018
rect 10222 5966 10274 6018
rect 12014 5966 12066 6018
rect 14478 5966 14530 6018
rect 7758 5854 7810 5906
rect 8094 5854 8146 5906
rect 12574 5854 12626 5906
rect 14590 5854 14642 5906
rect 2270 5742 2322 5794
rect 2718 5742 2770 5794
rect 8318 5742 8370 5794
rect 17614 5742 17666 5794
rect 18286 5742 18338 5794
rect 10446 5630 10498 5682
rect 3370 5462 3422 5514
rect 3474 5462 3526 5514
rect 3578 5462 3630 5514
rect 7682 5462 7734 5514
rect 7786 5462 7838 5514
rect 7890 5462 7942 5514
rect 11994 5462 12046 5514
rect 12098 5462 12150 5514
rect 12202 5462 12254 5514
rect 16306 5462 16358 5514
rect 16410 5462 16462 5514
rect 16514 5462 16566 5514
rect 11118 5294 11170 5346
rect 1710 5070 1762 5122
rect 3614 5070 3666 5122
rect 9550 5070 9602 5122
rect 10334 5070 10386 5122
rect 11006 5070 11058 5122
rect 16718 5070 16770 5122
rect 17166 5070 17218 5122
rect 18174 5070 18226 5122
rect 2046 4958 2098 5010
rect 9662 4958 9714 5010
rect 17838 4958 17890 5010
rect 2382 4846 2434 4898
rect 3166 4846 3218 4898
rect 15598 4846 15650 4898
rect 17614 4846 17666 4898
rect 5526 4678 5578 4730
rect 5630 4678 5682 4730
rect 5734 4678 5786 4730
rect 9838 4678 9890 4730
rect 9942 4678 9994 4730
rect 10046 4678 10098 4730
rect 14150 4678 14202 4730
rect 14254 4678 14306 4730
rect 14358 4678 14410 4730
rect 18462 4678 18514 4730
rect 18566 4678 18618 4730
rect 18670 4678 18722 4730
rect 2046 4510 2098 4562
rect 2718 4510 2770 4562
rect 5966 4510 6018 4562
rect 15710 4510 15762 4562
rect 16494 4510 16546 4562
rect 3054 4398 3106 4450
rect 17726 4398 17778 4450
rect 1710 4286 1762 4338
rect 2382 4286 2434 4338
rect 5630 4286 5682 4338
rect 15934 4286 15986 4338
rect 16830 4286 16882 4338
rect 17950 4286 18002 4338
rect 3838 4174 3890 4226
rect 4398 4174 4450 4226
rect 4846 4174 4898 4226
rect 5406 4174 5458 4226
rect 6414 4174 6466 4226
rect 6974 4174 7026 4226
rect 7646 4174 7698 4226
rect 8094 4174 8146 4226
rect 8654 4174 8706 4226
rect 9102 4174 9154 4226
rect 10110 4174 10162 4226
rect 10782 4174 10834 4226
rect 11454 4174 11506 4226
rect 13582 4174 13634 4226
rect 14254 4174 14306 4226
rect 14926 4174 14978 4226
rect 15486 4174 15538 4226
rect 3370 3894 3422 3946
rect 3474 3894 3526 3946
rect 3578 3894 3630 3946
rect 7682 3894 7734 3946
rect 7786 3894 7838 3946
rect 7890 3894 7942 3946
rect 11994 3894 12046 3946
rect 12098 3894 12150 3946
rect 12202 3894 12254 3946
rect 16306 3894 16358 3946
rect 16410 3894 16462 3946
rect 16514 3894 16566 3946
rect 1934 3502 1986 3554
rect 2718 3502 2770 3554
rect 3390 3502 3442 3554
rect 4062 3502 4114 3554
rect 4734 3502 4786 3554
rect 5854 3502 5906 3554
rect 6526 3502 6578 3554
rect 7198 3502 7250 3554
rect 7870 3502 7922 3554
rect 8654 3502 8706 3554
rect 9886 3502 9938 3554
rect 10558 3502 10610 3554
rect 11006 3502 11058 3554
rect 11902 3502 11954 3554
rect 12686 3502 12738 3554
rect 13358 3502 13410 3554
rect 14702 3502 14754 3554
rect 15486 3502 15538 3554
rect 16046 3502 16098 3554
rect 17166 3502 17218 3554
rect 2270 3390 2322 3442
rect 4958 3390 5010 3442
rect 8430 3390 8482 3442
rect 9662 3390 9714 3442
rect 11342 3390 11394 3442
rect 11678 3390 11730 3442
rect 13134 3390 13186 3442
rect 14142 3390 14194 3442
rect 14478 3390 14530 3442
rect 15150 3390 15202 3442
rect 15822 3390 15874 3442
rect 16942 3390 16994 3442
rect 17614 3390 17666 3442
rect 17950 3390 18002 3442
rect 2942 3278 2994 3330
rect 3614 3278 3666 3330
rect 4286 3278 4338 3330
rect 6078 3278 6130 3330
rect 6750 3278 6802 3330
rect 7422 3278 7474 3330
rect 8094 3278 8146 3330
rect 10334 3278 10386 3330
rect 13806 3278 13858 3330
rect 5526 3110 5578 3162
rect 5630 3110 5682 3162
rect 5734 3110 5786 3162
rect 9838 3110 9890 3162
rect 9942 3110 9994 3162
rect 10046 3110 10098 3162
rect 14150 3110 14202 3162
rect 14254 3110 14306 3162
rect 14358 3110 14410 3162
rect 18462 3110 18514 3162
rect 18566 3110 18618 3162
rect 18670 3110 18722 3162
rect 16830 2942 16882 2994
rect 17502 2942 17554 2994
rect 17950 2942 18002 2994
<< metal2 >>
rect 0 19200 112 20000
rect 672 19200 784 20000
rect 1344 19200 1456 20000
rect 2016 19200 2128 20000
rect 2688 19200 2800 20000
rect 3360 19200 3472 20000
rect 4032 19200 4144 20000
rect 4704 19200 4816 20000
rect 5376 19200 5488 20000
rect 6048 19200 6160 20000
rect 6720 19200 6832 20000
rect 7392 19200 7504 20000
rect 8064 19200 8176 20000
rect 8736 19200 8848 20000
rect 9408 19200 9520 20000
rect 10080 19200 10192 20000
rect 10752 19200 10864 20000
rect 11424 19200 11536 20000
rect 12096 19200 12208 20000
rect 12768 19200 12880 20000
rect 13440 19200 13552 20000
rect 14112 19200 14224 20000
rect 14784 19200 14896 20000
rect 15456 19200 15568 20000
rect 16128 19200 16240 20000
rect 16800 19200 16912 20000
rect 17472 19200 17584 20000
rect 18144 19200 18256 20000
rect 18816 19200 18928 20000
rect 19488 19200 19600 20000
rect 2716 16210 2772 19200
rect 3388 17332 3444 19200
rect 3388 17276 3780 17332
rect 3368 16492 3632 16502
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3368 16426 3632 16436
rect 2716 16158 2718 16210
rect 2770 16158 2772 16210
rect 2716 16146 2772 16158
rect 3164 16098 3220 16110
rect 3164 16046 3166 16098
rect 3218 16046 3220 16098
rect 1708 15876 1764 15886
rect 1708 15782 1764 15820
rect 1708 15426 1764 15438
rect 1708 15374 1710 15426
rect 1762 15374 1764 15426
rect 1708 15204 1764 15374
rect 1708 15138 1764 15148
rect 1708 14308 1764 14318
rect 1708 14214 1764 14252
rect 1708 13858 1764 13870
rect 1708 13806 1710 13858
rect 1762 13806 1764 13858
rect 1708 13524 1764 13806
rect 1708 13458 1764 13468
rect 1708 12290 1764 12302
rect 1708 12238 1710 12290
rect 1762 12238 1764 12290
rect 1708 11508 1764 12238
rect 1708 11442 1764 11452
rect 1820 11394 1876 11406
rect 1820 11342 1822 11394
rect 1874 11342 1876 11394
rect 1820 10836 1876 11342
rect 1820 10770 1876 10780
rect 2044 11170 2100 11182
rect 2044 11118 2046 11170
rect 2098 11118 2100 11170
rect 1708 10722 1764 10734
rect 1708 10670 1710 10722
rect 1762 10670 1764 10722
rect 1708 10164 1764 10670
rect 1708 10098 1764 10108
rect 2044 9828 2100 11118
rect 2492 11170 2548 11182
rect 2492 11118 2494 11170
rect 2546 11118 2548 11170
rect 2492 10836 2548 11118
rect 2492 10770 2548 10780
rect 3164 10052 3220 16046
rect 3612 15540 3668 15550
rect 3724 15540 3780 17276
rect 4060 16210 4116 19200
rect 4732 16324 4788 19200
rect 4732 16258 4788 16268
rect 4060 16158 4062 16210
rect 4114 16158 4116 16210
rect 4060 16146 4116 16158
rect 3612 15538 3780 15540
rect 3612 15486 3614 15538
rect 3666 15486 3780 15538
rect 3612 15484 3780 15486
rect 4956 16098 5012 16110
rect 4956 16046 4958 16098
rect 5010 16046 5012 16098
rect 3612 15474 3668 15484
rect 3368 14924 3632 14934
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3368 14858 3632 14868
rect 4956 13524 5012 16046
rect 5404 15540 5460 19200
rect 5964 16324 6020 16334
rect 5964 16230 6020 16268
rect 5524 15708 5788 15718
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5524 15642 5788 15652
rect 5628 15540 5684 15550
rect 5404 15538 5684 15540
rect 5404 15486 5630 15538
rect 5682 15486 5684 15538
rect 5404 15484 5684 15486
rect 6076 15540 6132 19200
rect 6748 17668 6804 19200
rect 6748 17612 7140 17668
rect 6636 16100 6692 16110
rect 6636 16006 6692 16044
rect 7084 15986 7140 17612
rect 7084 15934 7086 15986
rect 7138 15934 7140 15986
rect 7084 15922 7140 15934
rect 7420 16100 7476 19200
rect 7680 16492 7944 16502
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7680 16426 7944 16436
rect 7644 16100 7700 16110
rect 7420 16098 7700 16100
rect 7420 16046 7646 16098
rect 7698 16046 7700 16098
rect 7420 16044 7700 16046
rect 6300 15540 6356 15550
rect 6076 15538 6356 15540
rect 6076 15486 6302 15538
rect 6354 15486 6356 15538
rect 6076 15484 6356 15486
rect 5628 15474 5684 15484
rect 6300 15474 6356 15484
rect 7420 15538 7476 16044
rect 7644 16034 7700 16044
rect 7420 15486 7422 15538
rect 7474 15486 7476 15538
rect 7420 15474 7476 15486
rect 7980 15874 8036 15886
rect 7980 15822 7982 15874
rect 8034 15822 8036 15874
rect 7980 15148 8036 15822
rect 8092 15540 8148 19200
rect 8764 15986 8820 19200
rect 8764 15934 8766 15986
rect 8818 15934 8820 15986
rect 8764 15922 8820 15934
rect 9100 16100 9156 16110
rect 8316 15540 8372 15550
rect 8092 15538 8372 15540
rect 8092 15486 8318 15538
rect 8370 15486 8372 15538
rect 8092 15484 8372 15486
rect 8316 15474 8372 15484
rect 7980 15092 8148 15148
rect 7680 14924 7944 14934
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7680 14858 7944 14868
rect 6188 14418 6244 14430
rect 6188 14366 6190 14418
rect 6242 14366 6244 14418
rect 5524 14140 5788 14150
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5524 14074 5788 14084
rect 4956 13458 5012 13468
rect 3368 13356 3632 13366
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3368 13290 3632 13300
rect 5524 12572 5788 12582
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5524 12506 5788 12516
rect 4956 12180 5012 12190
rect 3368 11788 3632 11798
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3368 11722 3632 11732
rect 4956 11396 5012 12124
rect 6188 12178 6244 14366
rect 7680 13356 7944 13366
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7680 13290 7944 13300
rect 8092 12292 8148 15092
rect 8092 12226 8148 12236
rect 8988 13524 9044 13534
rect 6188 12126 6190 12178
rect 6242 12126 6244 12178
rect 6188 12114 6244 12126
rect 6076 12068 6132 12078
rect 5740 11956 5796 11966
rect 5740 11954 6020 11956
rect 5740 11902 5742 11954
rect 5794 11902 6020 11954
rect 5740 11900 6020 11902
rect 5740 11890 5796 11900
rect 5180 11396 5236 11406
rect 4956 11340 5180 11396
rect 5180 11302 5236 11340
rect 5740 11284 5796 11294
rect 5404 11282 5796 11284
rect 5404 11230 5742 11282
rect 5794 11230 5796 11282
rect 5404 11228 5796 11230
rect 5404 10836 5460 11228
rect 5740 11218 5796 11228
rect 5524 11004 5788 11014
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5524 10938 5788 10948
rect 5404 10780 5572 10836
rect 5404 10610 5460 10622
rect 5404 10558 5406 10610
rect 5458 10558 5460 10610
rect 3368 10220 3632 10230
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3368 10154 3632 10164
rect 3276 10052 3332 10062
rect 3164 9996 3276 10052
rect 3276 9986 3332 9996
rect 2044 9762 2100 9772
rect 5404 9044 5460 10558
rect 5516 10052 5572 10780
rect 5964 10610 6020 11900
rect 6076 11282 6132 12012
rect 6860 12068 6916 12078
rect 6860 11974 6916 12012
rect 8988 12066 9044 13468
rect 8988 12014 8990 12066
rect 9042 12014 9044 12066
rect 8316 11956 8372 11966
rect 7680 11788 7944 11798
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7680 11722 7944 11732
rect 6412 11396 6468 11406
rect 6412 11302 6468 11340
rect 6076 11230 6078 11282
rect 6130 11230 6132 11282
rect 6076 11218 6132 11230
rect 8316 10834 8372 11900
rect 8540 11172 8596 11182
rect 8316 10782 8318 10834
rect 8370 10782 8372 10834
rect 8316 10770 8372 10782
rect 8428 11116 8540 11172
rect 5964 10558 5966 10610
rect 6018 10558 6020 10610
rect 5964 10546 6020 10558
rect 5516 9986 5572 9996
rect 7532 10500 7588 10510
rect 8428 10500 8484 11116
rect 8540 11106 8596 11116
rect 8988 10612 9044 12014
rect 9100 10834 9156 16044
rect 9436 15988 9492 19200
rect 9660 15988 9716 15998
rect 9436 15986 9716 15988
rect 9436 15934 9662 15986
rect 9714 15934 9716 15986
rect 9436 15932 9716 15934
rect 10108 15988 10164 19200
rect 10780 16100 10836 19200
rect 11004 16100 11060 16110
rect 10780 16098 11060 16100
rect 10780 16046 11006 16098
rect 11058 16046 11060 16098
rect 10780 16044 11060 16046
rect 10332 15988 10388 15998
rect 10108 15986 10388 15988
rect 10108 15934 10334 15986
rect 10386 15934 10388 15986
rect 10108 15932 10388 15934
rect 9660 15922 9716 15932
rect 10332 15922 10388 15932
rect 9836 15708 10100 15718
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 9836 15642 10100 15652
rect 10780 15538 10836 16044
rect 11004 16034 11060 16044
rect 11452 15988 11508 19200
rect 12124 17556 12180 19200
rect 12796 17556 12852 19200
rect 12124 17500 12404 17556
rect 12796 17500 13188 17556
rect 11992 16492 12256 16502
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 11992 16426 12256 16436
rect 11676 15988 11732 15998
rect 11452 15986 11732 15988
rect 11452 15934 11678 15986
rect 11730 15934 11732 15986
rect 11452 15932 11732 15934
rect 11676 15922 11732 15932
rect 12348 15986 12404 17500
rect 12348 15934 12350 15986
rect 12402 15934 12404 15986
rect 12348 15922 12404 15934
rect 13132 15986 13188 17500
rect 13132 15934 13134 15986
rect 13186 15934 13188 15986
rect 13132 15922 13188 15934
rect 13468 15988 13524 19200
rect 13692 15988 13748 15998
rect 13468 15986 13748 15988
rect 13468 15934 13694 15986
rect 13746 15934 13748 15986
rect 13468 15932 13748 15934
rect 14140 15988 14196 19200
rect 14364 15988 14420 15998
rect 14140 15986 14420 15988
rect 14140 15934 14366 15986
rect 14418 15934 14420 15986
rect 14140 15932 14420 15934
rect 14812 15988 14868 19200
rect 15036 15988 15092 15998
rect 14812 15986 15092 15988
rect 14812 15934 15038 15986
rect 15090 15934 15092 15986
rect 14812 15932 15092 15934
rect 15484 15988 15540 19200
rect 15708 15988 15764 15998
rect 15484 15986 15764 15988
rect 15484 15934 15710 15986
rect 15762 15934 15764 15986
rect 15484 15932 15764 15934
rect 13692 15922 13748 15932
rect 14364 15922 14420 15932
rect 15036 15922 15092 15932
rect 15708 15922 15764 15932
rect 16156 15988 16212 19200
rect 16828 16770 16884 19200
rect 16828 16718 16830 16770
rect 16882 16718 16884 16770
rect 16828 16706 16884 16718
rect 17388 16770 17444 16782
rect 17388 16718 17390 16770
rect 17442 16718 17444 16770
rect 16304 16492 16568 16502
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16304 16426 16568 16436
rect 16156 15922 16212 15932
rect 16940 15988 16996 15998
rect 16940 15894 16996 15932
rect 17388 15986 17444 16718
rect 17388 15934 17390 15986
rect 17442 15934 17444 15986
rect 17388 15922 17444 15934
rect 17500 15988 17556 19200
rect 18172 17444 18228 19200
rect 17948 17388 18228 17444
rect 17836 15988 17892 15998
rect 17500 15986 17892 15988
rect 17500 15934 17838 15986
rect 17890 15934 17892 15986
rect 17500 15932 17892 15934
rect 17836 15922 17892 15932
rect 10780 15486 10782 15538
rect 10834 15486 10836 15538
rect 10780 15474 10836 15486
rect 11340 15874 11396 15886
rect 11340 15822 11342 15874
rect 11394 15822 11396 15874
rect 10444 14530 10500 14542
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 9836 14140 10100 14150
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 9836 14074 10100 14084
rect 9836 12572 10100 12582
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 9836 12506 10100 12516
rect 9884 12292 9940 12302
rect 9884 12198 9940 12236
rect 10332 12292 10388 12302
rect 10332 12198 10388 12236
rect 9772 11954 9828 11966
rect 9772 11902 9774 11954
rect 9826 11902 9828 11954
rect 9772 11172 9828 11902
rect 10220 11956 10276 11966
rect 10220 11862 10276 11900
rect 9772 11106 9828 11116
rect 10444 11282 10500 14478
rect 11340 11732 11396 15822
rect 16380 15876 16436 15886
rect 16380 15782 16436 15820
rect 17948 15764 18004 17388
rect 14148 15708 14412 15718
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14148 15642 14412 15652
rect 17724 15708 18004 15764
rect 18172 16770 18228 16782
rect 18172 16718 18174 16770
rect 18226 16718 18228 16770
rect 17724 15538 17780 15708
rect 17724 15486 17726 15538
rect 17778 15486 17780 15538
rect 17724 15474 17780 15486
rect 18172 15538 18228 16718
rect 18844 16770 18900 19200
rect 18844 16718 18846 16770
rect 18898 16718 18900 16770
rect 18844 16706 18900 16718
rect 19516 15876 19572 19200
rect 19516 15810 19572 15820
rect 18460 15708 18724 15718
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18460 15642 18724 15652
rect 18172 15486 18174 15538
rect 18226 15486 18228 15538
rect 18172 15474 18228 15486
rect 11992 14924 12256 14934
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 11992 14858 12256 14868
rect 16304 14924 16568 14934
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16304 14858 16568 14868
rect 14148 14140 14412 14150
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14148 14074 14412 14084
rect 18460 14140 18724 14150
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18460 14074 18724 14084
rect 11992 13356 12256 13366
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 11992 13290 12256 13300
rect 16304 13356 16568 13366
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16304 13290 16568 13300
rect 14148 12572 14412 12582
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14148 12506 14412 12516
rect 18460 12572 18724 12582
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18460 12506 18724 12516
rect 12236 12292 12292 12302
rect 12292 12236 12404 12292
rect 12236 12226 12292 12236
rect 11992 11788 12256 11798
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 11340 11676 11844 11732
rect 11992 11722 12256 11732
rect 10444 11230 10446 11282
rect 10498 11230 10500 11282
rect 9836 11004 10100 11014
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 9836 10938 10100 10948
rect 9100 10782 9102 10834
rect 9154 10782 9156 10834
rect 9100 10770 9156 10782
rect 9996 10722 10052 10734
rect 9996 10670 9998 10722
rect 10050 10670 10052 10722
rect 8988 10556 9604 10612
rect 7532 9828 7588 10444
rect 8316 10444 8484 10500
rect 7680 10220 7944 10230
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7680 10154 7944 10164
rect 7644 9828 7700 9838
rect 7532 9826 7700 9828
rect 7532 9774 7646 9826
rect 7698 9774 7700 9826
rect 7532 9772 7700 9774
rect 7644 9762 7700 9772
rect 8092 9826 8148 9838
rect 8092 9774 8094 9826
rect 8146 9774 8148 9826
rect 6076 9604 6132 9614
rect 5524 9436 5788 9446
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5524 9370 5788 9380
rect 5628 9044 5684 9054
rect 5404 9042 5684 9044
rect 5404 8990 5630 9042
rect 5682 8990 5684 9042
rect 5404 8988 5684 8990
rect 3368 8652 3632 8662
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3368 8586 3632 8596
rect 5628 8372 5684 8988
rect 6076 9042 6132 9548
rect 7420 9604 7476 9614
rect 7420 9510 7476 9548
rect 6076 8990 6078 9042
rect 6130 8990 6132 9042
rect 6076 8978 6132 8990
rect 7680 8652 7944 8662
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7680 8586 7944 8596
rect 5628 8306 5684 8316
rect 6636 8372 6692 8382
rect 6636 8278 6692 8316
rect 1708 8148 1764 8158
rect 1764 8092 1876 8148
rect 1708 8054 1764 8092
rect 1820 7698 1876 8092
rect 2044 8036 2100 8046
rect 2044 7942 2100 7980
rect 2380 8034 2436 8046
rect 2380 7982 2382 8034
rect 2434 7982 2436 8034
rect 1820 7646 1822 7698
rect 1874 7646 1876 7698
rect 1820 7634 1876 7646
rect 2380 7476 2436 7982
rect 5524 7868 5788 7878
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5524 7802 5788 7812
rect 7420 7586 7476 7598
rect 7420 7534 7422 7586
rect 7474 7534 7476 7586
rect 2380 7410 2436 7420
rect 2828 7476 2884 7486
rect 1820 6466 1876 6478
rect 1820 6414 1822 6466
rect 1874 6414 1876 6466
rect 1708 6018 1764 6030
rect 1708 5966 1710 6018
rect 1762 5966 1764 6018
rect 1708 5460 1764 5966
rect 1708 5394 1764 5404
rect 1708 5122 1764 5134
rect 1708 5070 1710 5122
rect 1762 5070 1764 5122
rect 812 5012 868 5022
rect 700 4956 812 5012
rect 28 3444 84 3454
rect 28 800 84 3388
rect 700 800 756 4956
rect 812 4946 868 4956
rect 1708 5012 1764 5070
rect 1708 4946 1764 4956
rect 1708 4340 1764 4350
rect 1820 4340 1876 6414
rect 2044 6468 2100 6478
rect 1708 4338 1876 4340
rect 1708 4286 1710 4338
rect 1762 4286 1876 4338
rect 1708 4284 1876 4286
rect 1932 5124 1988 5134
rect 1708 3668 1764 4284
rect 1372 3612 1764 3668
rect 1372 800 1428 3612
rect 1932 3556 1988 5068
rect 2044 5010 2100 6412
rect 2044 4958 2046 5010
rect 2098 4958 2100 5010
rect 2044 4946 2100 4958
rect 2268 5794 2324 5806
rect 2716 5796 2772 5806
rect 2268 5742 2270 5794
rect 2322 5742 2324 5794
rect 2268 5012 2324 5742
rect 2268 4946 2324 4956
rect 2604 5794 2772 5796
rect 2604 5742 2718 5794
rect 2770 5742 2772 5794
rect 2604 5740 2772 5742
rect 2380 4900 2436 4910
rect 2380 4806 2436 4844
rect 2044 4564 2100 4574
rect 2044 4470 2100 4508
rect 2268 4452 2324 4462
rect 1932 3554 2100 3556
rect 1932 3502 1934 3554
rect 1986 3502 2100 3554
rect 1932 3500 2100 3502
rect 1932 3490 1988 3500
rect 2044 800 2100 3500
rect 2268 3442 2324 4396
rect 2268 3390 2270 3442
rect 2322 3390 2324 3442
rect 2268 3378 2324 3390
rect 2380 4340 2436 4350
rect 2604 4340 2660 5740
rect 2716 5730 2772 5740
rect 2716 4564 2772 4574
rect 2828 4564 2884 7420
rect 7308 7474 7364 7486
rect 7308 7422 7310 7474
rect 7362 7422 7364 7474
rect 3368 7084 3632 7094
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3368 7018 3632 7028
rect 6748 6692 6804 6702
rect 2716 4562 2884 4564
rect 2716 4510 2718 4562
rect 2770 4510 2884 4562
rect 2716 4508 2884 4510
rect 2940 6580 2996 6590
rect 2716 4498 2772 4508
rect 2380 4338 2660 4340
rect 2380 4286 2382 4338
rect 2434 4286 2660 4338
rect 2380 4284 2660 4286
rect 2380 3444 2436 4284
rect 2380 3378 2436 3388
rect 2716 3554 2772 3566
rect 2716 3502 2718 3554
rect 2770 3502 2772 3554
rect 2716 3108 2772 3502
rect 2940 3330 2996 6524
rect 5524 6300 5788 6310
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5524 6234 5788 6244
rect 6076 6020 6132 6030
rect 3368 5516 3632 5526
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3368 5450 3632 5460
rect 3612 5124 3668 5134
rect 3612 5030 3668 5068
rect 4956 5012 5012 5022
rect 3164 4898 3220 4910
rect 3164 4846 3166 4898
rect 3218 4846 3220 4898
rect 3052 4450 3108 4462
rect 3052 4398 3054 4450
rect 3106 4398 3108 4450
rect 3052 4116 3108 4398
rect 3052 4050 3108 4060
rect 2940 3278 2942 3330
rect 2994 3278 2996 3330
rect 2940 3266 2996 3278
rect 3164 3108 3220 4846
rect 3836 4228 3892 4238
rect 4396 4228 4452 4238
rect 4844 4228 4900 4238
rect 3724 4226 3892 4228
rect 3724 4174 3838 4226
rect 3890 4174 3892 4226
rect 3724 4172 3892 4174
rect 3368 3948 3632 3958
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3368 3882 3632 3892
rect 3724 3668 3780 4172
rect 3836 4162 3892 4172
rect 4060 4226 4452 4228
rect 4060 4174 4398 4226
rect 4450 4174 4452 4226
rect 4060 4172 4452 4174
rect 2716 3052 3220 3108
rect 3388 3612 3780 3668
rect 3388 3554 3444 3612
rect 3388 3502 3390 3554
rect 3442 3502 3444 3554
rect 2716 800 2772 3052
rect 3388 800 3444 3502
rect 4060 3554 4116 4172
rect 4396 4162 4452 4172
rect 4732 4226 4900 4228
rect 4732 4174 4846 4226
rect 4898 4174 4900 4226
rect 4732 4172 4900 4174
rect 4060 3502 4062 3554
rect 4114 3502 4116 3554
rect 3612 3444 3668 3454
rect 3612 3330 3668 3388
rect 3612 3278 3614 3330
rect 3666 3278 3668 3330
rect 3612 3266 3668 3278
rect 4060 800 4116 3502
rect 4284 4004 4340 4014
rect 4284 3330 4340 3948
rect 4284 3278 4286 3330
rect 4338 3278 4340 3330
rect 4284 3266 4340 3278
rect 4732 3554 4788 4172
rect 4844 4162 4900 4172
rect 4732 3502 4734 3554
rect 4786 3502 4788 3554
rect 4732 800 4788 3502
rect 4956 3442 5012 4956
rect 5964 4900 6020 4910
rect 5524 4732 5788 4742
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5524 4666 5788 4676
rect 5964 4562 6020 4844
rect 5964 4510 5966 4562
rect 6018 4510 6020 4562
rect 5964 4498 6020 4510
rect 5628 4338 5684 4350
rect 5628 4286 5630 4338
rect 5682 4286 5684 4338
rect 4956 3390 4958 3442
rect 5010 3390 5012 3442
rect 4956 3378 5012 3390
rect 5404 4228 5460 4238
rect 5628 4228 5684 4286
rect 5404 4226 5684 4228
rect 5404 4174 5406 4226
rect 5458 4174 5684 4226
rect 5404 4172 5684 4174
rect 5404 800 5460 4172
rect 5852 3554 5908 3566
rect 5852 3502 5854 3554
rect 5906 3502 5908 3554
rect 5524 3164 5788 3174
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5524 3098 5788 3108
rect 5852 3108 5908 3502
rect 6076 3330 6132 5964
rect 6412 4228 6468 4238
rect 6300 4226 6468 4228
rect 6300 4174 6414 4226
rect 6466 4174 6468 4226
rect 6300 4172 6468 4174
rect 6300 3388 6356 4172
rect 6412 4162 6468 4172
rect 6524 3554 6580 3566
rect 6524 3502 6526 3554
rect 6578 3502 6580 3554
rect 6524 3388 6580 3502
rect 6300 3332 6468 3388
rect 6524 3332 6692 3388
rect 6076 3278 6078 3330
rect 6130 3278 6132 3330
rect 6076 3266 6132 3278
rect 6412 3108 6468 3332
rect 5852 3052 6468 3108
rect 6636 3108 6692 3332
rect 6748 3330 6804 6636
rect 7084 6020 7140 6030
rect 7084 5926 7140 5964
rect 7308 4564 7364 7422
rect 7420 6468 7476 7534
rect 8092 7252 8148 9774
rect 7420 6402 7476 6412
rect 7532 7196 8148 7252
rect 8204 9714 8260 9726
rect 8204 9662 8206 9714
rect 8258 9662 8260 9714
rect 7532 5124 7588 7196
rect 7680 7084 7944 7094
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7680 7018 7944 7028
rect 8204 6916 8260 9662
rect 8316 9266 8372 10444
rect 8316 9214 8318 9266
rect 8370 9214 8372 9266
rect 8316 9202 8372 9214
rect 9100 9940 9156 9950
rect 9100 9268 9156 9884
rect 9100 9174 9156 9212
rect 9548 9044 9604 10556
rect 9884 10610 9940 10622
rect 9884 10558 9886 10610
rect 9938 10558 9940 10610
rect 9660 10052 9716 10062
rect 9660 9266 9716 9996
rect 9884 9604 9940 10558
rect 9996 10612 10052 10670
rect 9996 10556 10164 10612
rect 9996 10388 10052 10398
rect 9996 10294 10052 10332
rect 10108 9604 10164 10556
rect 10332 10276 10388 10286
rect 10108 9548 10276 9604
rect 9884 9538 9940 9548
rect 9836 9436 10100 9446
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 9836 9370 10100 9380
rect 9660 9214 9662 9266
rect 9714 9214 9716 9266
rect 9660 9202 9716 9214
rect 9996 9044 10052 9054
rect 9548 9042 10052 9044
rect 9548 8990 9998 9042
rect 10050 8990 10052 9042
rect 9548 8988 10052 8990
rect 9996 8978 10052 8988
rect 9836 7868 10100 7878
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 9836 7802 10100 7812
rect 10220 7700 10276 9548
rect 10332 9154 10388 10220
rect 10332 9102 10334 9154
rect 10386 9102 10388 9154
rect 10332 9090 10388 9102
rect 10444 8258 10500 11230
rect 11788 10722 11844 11676
rect 11788 10670 11790 10722
rect 11842 10670 11844 10722
rect 11788 10658 11844 10670
rect 11676 10610 11732 10622
rect 11676 10558 11678 10610
rect 11730 10558 11732 10610
rect 10892 10500 10948 10510
rect 10892 10406 10948 10444
rect 10556 10388 10612 10398
rect 10556 9492 10612 10332
rect 11228 10386 11284 10398
rect 11228 10334 11230 10386
rect 11282 10334 11284 10386
rect 10668 9714 10724 9726
rect 10668 9662 10670 9714
rect 10722 9662 10724 9714
rect 10668 9604 10724 9662
rect 10668 9548 10836 9604
rect 10556 9436 10724 9492
rect 10556 9268 10612 9278
rect 10556 9154 10612 9212
rect 10556 9102 10558 9154
rect 10610 9102 10612 9154
rect 10556 9090 10612 9102
rect 10444 8206 10446 8258
rect 10498 8206 10500 8258
rect 10444 8194 10500 8206
rect 10108 7644 10276 7700
rect 8988 7586 9044 7598
rect 8988 7534 8990 7586
rect 9042 7534 9044 7586
rect 8428 7476 8484 7486
rect 8428 7382 8484 7420
rect 8092 6860 8260 6916
rect 8316 7362 8372 7374
rect 8316 7310 8318 7362
rect 8370 7310 8372 7362
rect 8092 6132 8148 6860
rect 8316 6804 8372 7310
rect 8316 6748 8484 6804
rect 8204 6692 8260 6702
rect 8204 6598 8260 6636
rect 8092 6076 8260 6132
rect 7756 5906 7812 5918
rect 7756 5854 7758 5906
rect 7810 5854 7812 5906
rect 7756 5684 7812 5854
rect 8092 5908 8148 5918
rect 8092 5814 8148 5852
rect 7756 5628 8148 5684
rect 7680 5516 7944 5526
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7680 5450 7944 5460
rect 7308 4498 7364 4508
rect 7420 5068 7588 5124
rect 6748 3278 6750 3330
rect 6802 3278 6804 3330
rect 6748 3266 6804 3278
rect 6972 4226 7028 4238
rect 6972 4174 6974 4226
rect 7026 4174 7028 4226
rect 6972 3108 7028 4174
rect 6636 3052 7028 3108
rect 7196 3554 7252 3566
rect 7196 3502 7198 3554
rect 7250 3502 7252 3554
rect 7196 3108 7252 3502
rect 7420 3330 7476 5068
rect 8092 4676 8148 5628
rect 8092 4610 8148 4620
rect 7644 4228 7700 4238
rect 7420 3278 7422 3330
rect 7474 3278 7476 3330
rect 7420 3266 7476 3278
rect 7532 4226 7700 4228
rect 7532 4174 7646 4226
rect 7698 4174 7700 4226
rect 7532 4172 7700 4174
rect 7532 3108 7588 4172
rect 7644 4162 7700 4172
rect 8092 4226 8148 4238
rect 8092 4174 8094 4226
rect 8146 4174 8148 4226
rect 7680 3948 7944 3958
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7680 3882 7944 3892
rect 7196 3052 7588 3108
rect 5852 2324 5908 3052
rect 5852 2268 6132 2324
rect 6076 800 6132 2268
rect 6748 800 6804 3052
rect 7532 2548 7588 3052
rect 7420 2492 7588 2548
rect 7868 3556 7924 3566
rect 8092 3556 8148 4174
rect 7868 3554 8148 3556
rect 7868 3502 7870 3554
rect 7922 3502 8148 3554
rect 7868 3500 8148 3502
rect 7420 800 7476 2492
rect 7868 980 7924 3500
rect 8204 3388 8260 6076
rect 8316 5796 8372 5806
rect 8316 5702 8372 5740
rect 8428 5124 8484 6748
rect 8764 6580 8820 6590
rect 8652 6578 8820 6580
rect 8652 6526 8766 6578
rect 8818 6526 8820 6578
rect 8652 6524 8820 6526
rect 8428 5058 8484 5068
rect 8540 5908 8596 5918
rect 8092 3332 8260 3388
rect 8428 4676 8484 4686
rect 8428 3442 8484 4620
rect 8540 4452 8596 5852
rect 8652 5012 8708 6524
rect 8764 6514 8820 6524
rect 8764 6020 8820 6030
rect 8764 6018 8932 6020
rect 8764 5966 8766 6018
rect 8818 5966 8932 6018
rect 8764 5964 8932 5966
rect 8764 5954 8820 5964
rect 8652 4946 8708 4956
rect 8540 4386 8596 4396
rect 8428 3390 8430 3442
rect 8482 3390 8484 3442
rect 8428 3378 8484 3390
rect 8652 4226 8708 4238
rect 8652 4174 8654 4226
rect 8706 4174 8708 4226
rect 8652 3554 8708 4174
rect 8652 3502 8654 3554
rect 8706 3502 8708 3554
rect 8652 3388 8708 3502
rect 8876 3444 8932 5964
rect 8988 5460 9044 7534
rect 9884 7476 9940 7486
rect 8988 5394 9044 5404
rect 9436 7474 9940 7476
rect 9436 7422 9886 7474
rect 9938 7422 9940 7474
rect 9436 7420 9940 7422
rect 9100 4228 9156 4238
rect 9100 4134 9156 4172
rect 9436 3780 9492 7420
rect 9884 7410 9940 7420
rect 9996 7362 10052 7374
rect 9996 7310 9998 7362
rect 10050 7310 10052 7362
rect 9996 6692 10052 7310
rect 10108 7028 10164 7644
rect 10556 7476 10612 7486
rect 10668 7476 10724 9436
rect 10556 7474 10724 7476
rect 10556 7422 10558 7474
rect 10610 7422 10724 7474
rect 10556 7420 10724 7422
rect 10556 7410 10612 7420
rect 10220 7250 10276 7262
rect 10220 7198 10222 7250
rect 10274 7198 10276 7250
rect 10220 7140 10276 7198
rect 10220 7084 10612 7140
rect 10108 6972 10388 7028
rect 9996 6626 10052 6636
rect 10220 6690 10276 6702
rect 10220 6638 10222 6690
rect 10274 6638 10276 6690
rect 9660 6466 9716 6478
rect 9660 6414 9662 6466
rect 9714 6414 9716 6466
rect 9548 5124 9604 5134
rect 9548 5030 9604 5068
rect 9660 5010 9716 6414
rect 9836 6300 10100 6310
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 9836 6234 10100 6244
rect 10220 6244 10276 6638
rect 10220 6178 10276 6188
rect 10332 6130 10388 6972
rect 10332 6078 10334 6130
rect 10386 6078 10388 6130
rect 10332 6066 10388 6078
rect 9660 4958 9662 5010
rect 9714 4958 9716 5010
rect 9660 4946 9716 4958
rect 10220 6018 10276 6030
rect 10220 5966 10222 6018
rect 10274 5966 10276 6018
rect 9836 4732 10100 4742
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 9836 4666 10100 4676
rect 10220 4452 10276 5966
rect 10332 5796 10388 5806
rect 10332 5122 10388 5740
rect 10444 5684 10500 5694
rect 10444 5590 10500 5628
rect 10332 5070 10334 5122
rect 10386 5070 10388 5122
rect 10332 5058 10388 5070
rect 10444 5460 10500 5470
rect 10220 4386 10276 4396
rect 9436 3714 9492 3724
rect 9884 4228 9940 4238
rect 9884 3554 9940 4172
rect 9884 3502 9886 3554
rect 9938 3502 9940 3554
rect 9660 3444 9716 3454
rect 8876 3442 9716 3444
rect 8876 3390 9662 3442
rect 9714 3390 9716 3442
rect 8876 3388 9716 3390
rect 8652 3332 8820 3388
rect 9660 3378 9716 3388
rect 8092 3330 8148 3332
rect 8092 3278 8094 3330
rect 8146 3278 8148 3330
rect 8092 3266 8148 3278
rect 7868 924 8148 980
rect 8092 800 8148 924
rect 8764 800 8820 3332
rect 9884 3332 9940 3502
rect 10108 4226 10164 4238
rect 10108 4174 10110 4226
rect 10162 4174 10164 4226
rect 10108 3388 10164 4174
rect 10444 3388 10500 5404
rect 10556 4228 10612 7084
rect 10780 6804 10836 9548
rect 11116 9602 11172 9614
rect 11116 9550 11118 9602
rect 11170 9550 11172 9602
rect 11116 7812 11172 9550
rect 11228 9268 11284 10334
rect 11676 10052 11732 10558
rect 11992 10220 12256 10230
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 11992 10154 12256 10164
rect 11676 9986 11732 9996
rect 12236 10052 12292 10062
rect 12348 10052 12404 12236
rect 16304 11788 16568 11798
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16304 11722 16568 11732
rect 14148 11004 14412 11014
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14148 10938 14412 10948
rect 18460 11004 18724 11014
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18460 10938 18724 10948
rect 12572 10724 12628 10734
rect 12572 10722 12740 10724
rect 12572 10670 12574 10722
rect 12626 10670 12740 10722
rect 12572 10668 12740 10670
rect 12572 10658 12628 10668
rect 12236 10050 12404 10052
rect 12236 9998 12238 10050
rect 12290 9998 12404 10050
rect 12236 9996 12404 9998
rect 12460 10610 12516 10622
rect 12460 10558 12462 10610
rect 12514 10558 12516 10610
rect 12236 9986 12292 9996
rect 12460 9938 12516 10558
rect 12572 10388 12628 10398
rect 12572 10294 12628 10332
rect 12460 9886 12462 9938
rect 12514 9886 12516 9938
rect 12460 9874 12516 9886
rect 11900 9828 11956 9838
rect 11228 9202 11284 9212
rect 11564 9826 11956 9828
rect 11564 9774 11902 9826
rect 11954 9774 11956 9826
rect 11564 9772 11956 9774
rect 12684 9828 12740 10668
rect 16304 10220 16568 10230
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16304 10154 16568 10164
rect 13468 10052 13524 10062
rect 12796 9828 12852 9838
rect 12684 9772 12796 9828
rect 10668 6748 10836 6804
rect 11004 7756 11172 7812
rect 11340 9154 11396 9166
rect 11340 9102 11342 9154
rect 11394 9102 11396 9154
rect 10668 6356 10724 6748
rect 10780 6580 10836 6590
rect 10780 6486 10836 6524
rect 10668 6300 10836 6356
rect 10556 4162 10612 4172
rect 10668 6132 10724 6142
rect 10108 3332 10276 3388
rect 9884 3266 9940 3276
rect 9436 3220 9492 3230
rect 9436 800 9492 3164
rect 9836 3164 10100 3174
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 9836 3098 10100 3108
rect 10220 3108 10276 3332
rect 10332 3332 10500 3388
rect 10556 3554 10612 3566
rect 10556 3502 10558 3554
rect 10610 3502 10612 3554
rect 10332 3330 10388 3332
rect 10332 3278 10334 3330
rect 10386 3278 10388 3330
rect 10332 3266 10388 3278
rect 10556 3108 10612 3502
rect 10668 3444 10724 6076
rect 10780 4452 10836 6300
rect 11004 5122 11060 7756
rect 11116 7586 11172 7598
rect 11116 7534 11118 7586
rect 11170 7534 11172 7586
rect 11116 5346 11172 7534
rect 11116 5294 11118 5346
rect 11170 5294 11172 5346
rect 11116 5282 11172 5294
rect 11004 5070 11006 5122
rect 11058 5070 11060 5122
rect 11004 5058 11060 5070
rect 10780 4396 10948 4452
rect 10668 3378 10724 3388
rect 10780 4226 10836 4238
rect 10780 4174 10782 4226
rect 10834 4174 10836 4226
rect 10780 3556 10836 4174
rect 10892 4116 10948 4396
rect 10892 4050 10948 4060
rect 11004 3556 11060 3566
rect 10780 3554 11060 3556
rect 10780 3502 11006 3554
rect 11058 3502 11060 3554
rect 10780 3500 11060 3502
rect 10220 3052 10612 3108
rect 10220 2884 10276 3052
rect 10108 2828 10276 2884
rect 10108 800 10164 2828
rect 10780 800 10836 3500
rect 11004 3490 11060 3500
rect 11340 3442 11396 9102
rect 11564 4900 11620 9772
rect 11900 9762 11956 9772
rect 12796 9762 12852 9772
rect 13356 9828 13412 9838
rect 13468 9828 13524 9996
rect 13356 9826 13524 9828
rect 13356 9774 13358 9826
rect 13410 9774 13524 9826
rect 13356 9772 13524 9774
rect 13692 9828 13748 9838
rect 13356 9762 13412 9772
rect 12460 9716 12516 9726
rect 12460 9622 12516 9660
rect 13580 9716 13636 9726
rect 13580 9622 13636 9660
rect 13692 9716 13748 9772
rect 13692 9714 13860 9716
rect 13692 9662 13694 9714
rect 13746 9662 13860 9714
rect 13692 9660 13860 9662
rect 13692 9650 13748 9660
rect 11788 9604 11844 9614
rect 11788 9266 11844 9548
rect 11788 9214 11790 9266
rect 11842 9214 11844 9266
rect 11788 9202 11844 9214
rect 12684 9156 12740 9166
rect 11788 9044 11844 9054
rect 11564 4834 11620 4844
rect 11676 9042 11844 9044
rect 11676 8990 11790 9042
rect 11842 8990 11844 9042
rect 11676 8988 11844 8990
rect 11340 3390 11342 3442
rect 11394 3390 11396 3442
rect 11340 3378 11396 3390
rect 11452 4226 11508 4238
rect 11452 4174 11454 4226
rect 11506 4174 11508 4226
rect 11452 3556 11508 4174
rect 11452 800 11508 3500
rect 11676 3442 11732 8988
rect 11788 8978 11844 8988
rect 12348 9042 12404 9054
rect 12348 8990 12350 9042
rect 12402 8990 12404 9042
rect 11992 8652 12256 8662
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 11992 8586 12256 8596
rect 11992 7084 12256 7094
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 11992 7018 12256 7028
rect 12012 6020 12068 6030
rect 12012 5926 12068 5964
rect 11992 5516 12256 5526
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 11992 5450 12256 5460
rect 12348 5012 12404 8990
rect 12684 8370 12740 9100
rect 12684 8318 12686 8370
rect 12738 8318 12740 8370
rect 12684 8306 12740 8318
rect 12796 9154 12852 9166
rect 12796 9102 12798 9154
rect 12850 9102 12852 9154
rect 12572 8260 12628 8270
rect 12460 8258 12628 8260
rect 12460 8206 12574 8258
rect 12626 8206 12628 8258
rect 12460 8204 12628 8206
rect 12460 5572 12516 8204
rect 12572 8194 12628 8204
rect 12684 8036 12740 8046
rect 12572 6692 12628 6702
rect 12572 6598 12628 6636
rect 12684 6578 12740 7980
rect 12684 6526 12686 6578
rect 12738 6526 12740 6578
rect 12684 6514 12740 6526
rect 12796 6356 12852 9102
rect 13468 9156 13524 9166
rect 13468 9062 13524 9100
rect 13356 9042 13412 9054
rect 13356 8990 13358 9042
rect 13410 8990 13412 9042
rect 13356 8932 13412 8990
rect 13356 8876 13524 8932
rect 12908 8148 12964 8158
rect 12908 8146 13412 8148
rect 12908 8094 12910 8146
rect 12962 8094 13412 8146
rect 12908 8092 13412 8094
rect 12908 8082 12964 8092
rect 13132 7586 13188 7598
rect 13132 7534 13134 7586
rect 13186 7534 13188 7586
rect 13132 6804 13188 7534
rect 12908 6748 13188 6804
rect 12908 6690 12964 6748
rect 12908 6638 12910 6690
rect 12962 6638 12964 6690
rect 12908 6626 12964 6638
rect 12796 6300 13188 6356
rect 12572 5908 12628 5918
rect 12572 5814 12628 5852
rect 12460 5506 12516 5516
rect 12460 5012 12516 5022
rect 12348 4956 12460 5012
rect 12460 4946 12516 4956
rect 11992 3948 12256 3958
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 11992 3882 12256 3892
rect 11900 3556 11956 3566
rect 11900 3462 11956 3500
rect 12684 3556 12740 3566
rect 11676 3390 11678 3442
rect 11730 3390 11732 3442
rect 11676 3378 11732 3390
rect 12684 3388 12740 3500
rect 12124 3332 12740 3388
rect 12796 3444 12852 3454
rect 12124 800 12180 3332
rect 12796 800 12852 3388
rect 13132 3442 13188 6300
rect 13356 5796 13412 8092
rect 13468 7476 13524 8876
rect 13804 7698 13860 9660
rect 14148 9436 14412 9446
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14148 9370 14412 9380
rect 18460 9436 18724 9446
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18460 9370 18724 9380
rect 17836 9154 17892 9166
rect 17836 9102 17838 9154
rect 17890 9102 17892 9154
rect 13916 9042 13972 9054
rect 13916 8990 13918 9042
rect 13970 8990 13972 9042
rect 13916 8260 13972 8990
rect 14700 9042 14756 9054
rect 14700 8990 14702 9042
rect 14754 8990 14756 9042
rect 13916 8194 13972 8204
rect 14476 8818 14532 8830
rect 14476 8766 14478 8818
rect 14530 8766 14532 8818
rect 14148 7868 14412 7878
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14148 7802 14412 7812
rect 13804 7646 13806 7698
rect 13858 7646 13860 7698
rect 13804 7634 13860 7646
rect 14364 7476 14420 7486
rect 14476 7476 14532 8766
rect 14700 8148 14756 8990
rect 17612 8930 17668 8942
rect 17612 8878 17614 8930
rect 17666 8878 17668 8930
rect 17612 8820 17668 8878
rect 17612 8754 17668 8764
rect 16304 8652 16568 8662
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16304 8586 16568 8596
rect 17836 8428 17892 9102
rect 18172 9042 18228 9054
rect 18172 8990 18174 9042
rect 18226 8990 18228 9042
rect 18172 8820 18228 8990
rect 18172 8754 18228 8764
rect 17836 8372 18004 8428
rect 14700 8082 14756 8092
rect 17164 8260 17220 8270
rect 17164 8146 17220 8204
rect 17164 8094 17166 8146
rect 17218 8094 17220 8146
rect 17164 8082 17220 8094
rect 17500 8146 17556 8158
rect 17500 8094 17502 8146
rect 17554 8094 17556 8146
rect 13468 7420 13636 7476
rect 13580 6130 13636 7420
rect 14364 7474 14532 7476
rect 14364 7422 14366 7474
rect 14418 7422 14532 7474
rect 14364 7420 14532 7422
rect 17500 7476 17556 8094
rect 17836 8148 17892 8158
rect 17836 8054 17892 8092
rect 17724 7476 17780 7486
rect 17500 7420 17724 7476
rect 14364 7410 14420 7420
rect 17724 7382 17780 7420
rect 16304 7084 16568 7094
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16304 7018 16568 7028
rect 14148 6300 14412 6310
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14148 6234 14412 6244
rect 13580 6078 13582 6130
rect 13634 6078 13636 6130
rect 13580 6066 13636 6078
rect 14476 6018 14532 6030
rect 14476 5966 14478 6018
rect 14530 5966 14532 6018
rect 13356 5740 13860 5796
rect 13580 4226 13636 4238
rect 13580 4174 13582 4226
rect 13634 4174 13636 4226
rect 13356 3556 13412 3566
rect 13356 3462 13412 3500
rect 13132 3390 13134 3442
rect 13186 3390 13188 3442
rect 13132 3378 13188 3390
rect 13580 3444 13636 4174
rect 13580 3378 13636 3388
rect 13804 3330 13860 5740
rect 14148 4732 14412 4742
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14148 4666 14412 4676
rect 14252 4228 14308 4238
rect 13804 3278 13806 3330
rect 13858 3278 13860 3330
rect 13804 3266 13860 3278
rect 14028 4226 14308 4228
rect 14028 4174 14254 4226
rect 14306 4174 14308 4226
rect 14028 4172 14308 4174
rect 14028 2996 14084 4172
rect 14252 4162 14308 4172
rect 14140 3444 14196 3482
rect 14140 3378 14196 3388
rect 14476 3442 14532 5966
rect 17948 6020 18004 8372
rect 18172 8148 18228 8158
rect 18228 8092 18340 8148
rect 18172 8054 18228 8092
rect 18284 7698 18340 8092
rect 18460 7868 18724 7878
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18460 7802 18724 7812
rect 18284 7646 18286 7698
rect 18338 7646 18340 7698
rect 18284 7634 18340 7646
rect 18460 6300 18724 6310
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18460 6234 18724 6244
rect 17948 5954 18004 5964
rect 14588 5906 14644 5918
rect 14588 5854 14590 5906
rect 14642 5854 14644 5906
rect 14588 4564 14644 5854
rect 14588 4498 14644 4508
rect 15148 5908 15204 5918
rect 14924 4228 14980 4238
rect 14812 4226 14980 4228
rect 14812 4174 14926 4226
rect 14978 4174 14980 4226
rect 14812 4172 14980 4174
rect 14476 3390 14478 3442
rect 14530 3390 14532 3442
rect 14476 3378 14532 3390
rect 14700 3554 14756 3566
rect 14700 3502 14702 3554
rect 14754 3502 14756 3554
rect 14148 3164 14412 3174
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14148 3098 14412 3108
rect 14700 2996 14756 3502
rect 14028 2940 14756 2996
rect 14812 3556 14868 4172
rect 14924 4162 14980 4172
rect 14028 2324 14084 2940
rect 13468 2268 14084 2324
rect 13468 800 13524 2268
rect 14812 1876 14868 3500
rect 14140 1820 14868 1876
rect 14924 3444 14980 3454
rect 14140 800 14196 1820
rect 14924 1764 14980 3388
rect 15148 3442 15204 5852
rect 17612 5796 17668 5806
rect 17500 5794 17668 5796
rect 17500 5742 17614 5794
rect 17666 5742 17668 5794
rect 17500 5740 17668 5742
rect 16044 5572 16100 5582
rect 15596 4900 15652 4910
rect 15148 3390 15150 3442
rect 15202 3390 15204 3442
rect 15148 3378 15204 3390
rect 15372 4898 15652 4900
rect 15372 4846 15598 4898
rect 15650 4846 15652 4898
rect 15372 4844 15652 4846
rect 15372 3444 15428 4844
rect 15596 4834 15652 4844
rect 15708 4564 15764 4574
rect 15708 4470 15764 4508
rect 15932 4338 15988 4350
rect 15932 4286 15934 4338
rect 15986 4286 15988 4338
rect 15484 4228 15540 4238
rect 15932 4228 15988 4286
rect 15484 4226 15988 4228
rect 15484 4174 15486 4226
rect 15538 4174 15988 4226
rect 15484 4172 15988 4174
rect 15484 4162 15540 4172
rect 15484 3556 15540 3566
rect 15484 3462 15540 3500
rect 15372 3378 15428 3388
rect 15596 3332 15652 4172
rect 16044 4116 16100 5516
rect 16304 5516 16568 5526
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16304 5450 16568 5460
rect 16716 5122 16772 5134
rect 16716 5070 16718 5122
rect 16770 5070 16772 5122
rect 16492 5012 16548 5022
rect 16492 4562 16548 4956
rect 16492 4510 16494 4562
rect 16546 4510 16548 4562
rect 16492 4498 16548 4510
rect 15820 4060 16100 4116
rect 15820 3442 15876 4060
rect 16304 3948 16568 3958
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16304 3882 16568 3892
rect 15820 3390 15822 3442
rect 15874 3390 15876 3442
rect 15820 3378 15876 3390
rect 16044 3554 16100 3566
rect 16044 3502 16046 3554
rect 16098 3502 16100 3554
rect 16044 3444 16100 3502
rect 16044 3378 16100 3388
rect 16268 3444 16324 3454
rect 14812 1708 14980 1764
rect 15484 3276 15652 3332
rect 14812 800 14868 1708
rect 15484 800 15540 3276
rect 16268 3220 16324 3388
rect 16716 3444 16772 5070
rect 17164 5122 17220 5134
rect 17164 5070 17166 5122
rect 17218 5070 17220 5122
rect 16828 4340 16884 4350
rect 16828 4246 16884 4284
rect 17164 4340 17220 5070
rect 17164 4274 17220 4284
rect 16716 3378 16772 3388
rect 16940 3780 16996 3790
rect 16940 3442 16996 3724
rect 16940 3390 16942 3442
rect 16994 3390 16996 3442
rect 16940 3378 16996 3390
rect 17164 3554 17220 3566
rect 17164 3502 17166 3554
rect 17218 3502 17220 3554
rect 17164 3444 17220 3502
rect 17164 3378 17220 3388
rect 16156 3164 16324 3220
rect 16156 800 16212 3164
rect 16828 2994 16884 3006
rect 16828 2942 16830 2994
rect 16882 2942 16884 2994
rect 16828 800 16884 2942
rect 17500 2994 17556 5740
rect 17612 5730 17668 5740
rect 18284 5794 18340 5806
rect 18284 5742 18286 5794
rect 18338 5742 18340 5794
rect 17836 5684 17892 5694
rect 17836 5010 17892 5628
rect 17836 4958 17838 5010
rect 17890 4958 17892 5010
rect 17836 4946 17892 4958
rect 18172 5124 18228 5134
rect 18284 5124 18340 5742
rect 18172 5122 18340 5124
rect 18172 5070 18174 5122
rect 18226 5070 18340 5122
rect 18172 5068 18340 5070
rect 17612 4898 17668 4910
rect 17612 4846 17614 4898
rect 17666 4846 17668 4898
rect 17612 4676 17668 4846
rect 17612 4620 17892 4676
rect 17724 4452 17780 4462
rect 17724 4358 17780 4396
rect 17836 4340 17892 4620
rect 17948 4340 18004 4350
rect 17836 4338 18004 4340
rect 17836 4286 17950 4338
rect 18002 4286 18004 4338
rect 17836 4284 18004 4286
rect 17612 4228 17668 4238
rect 17612 3442 17668 4172
rect 17612 3390 17614 3442
rect 17666 3390 17668 3442
rect 17612 3378 17668 3390
rect 17500 2942 17502 2994
rect 17554 2942 17556 2994
rect 17500 2930 17556 2942
rect 17836 2772 17892 4284
rect 17948 4274 18004 4284
rect 18060 4340 18116 4350
rect 17948 3442 18004 3454
rect 17948 3390 17950 3442
rect 18002 3390 18004 3442
rect 17948 2994 18004 3390
rect 17948 2942 17950 2994
rect 18002 2942 18004 2994
rect 17948 2930 18004 2942
rect 18060 2884 18116 4284
rect 18172 3668 18228 5068
rect 18460 4732 18724 4742
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18460 4666 18724 4676
rect 18172 3612 18900 3668
rect 18460 3164 18724 3174
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18460 3098 18724 3108
rect 18060 2828 18228 2884
rect 17500 2716 17892 2772
rect 17500 800 17556 2716
rect 18172 800 18228 2828
rect 18844 800 18900 3612
rect 0 0 112 800
rect 672 0 784 800
rect 1344 0 1456 800
rect 2016 0 2128 800
rect 2688 0 2800 800
rect 3360 0 3472 800
rect 4032 0 4144 800
rect 4704 0 4816 800
rect 5376 0 5488 800
rect 6048 0 6160 800
rect 6720 0 6832 800
rect 7392 0 7504 800
rect 8064 0 8176 800
rect 8736 0 8848 800
rect 9408 0 9520 800
rect 10080 0 10192 800
rect 10752 0 10864 800
rect 11424 0 11536 800
rect 12096 0 12208 800
rect 12768 0 12880 800
rect 13440 0 13552 800
rect 14112 0 14224 800
rect 14784 0 14896 800
rect 15456 0 15568 800
rect 16128 0 16240 800
rect 16800 0 16912 800
rect 17472 0 17584 800
rect 18144 0 18256 800
rect 18816 0 18928 800
rect 19488 0 19600 800
<< via2 >>
rect 3368 16490 3424 16492
rect 3368 16438 3370 16490
rect 3370 16438 3422 16490
rect 3422 16438 3424 16490
rect 3368 16436 3424 16438
rect 3472 16490 3528 16492
rect 3472 16438 3474 16490
rect 3474 16438 3526 16490
rect 3526 16438 3528 16490
rect 3472 16436 3528 16438
rect 3576 16490 3632 16492
rect 3576 16438 3578 16490
rect 3578 16438 3630 16490
rect 3630 16438 3632 16490
rect 3576 16436 3632 16438
rect 1708 15874 1764 15876
rect 1708 15822 1710 15874
rect 1710 15822 1762 15874
rect 1762 15822 1764 15874
rect 1708 15820 1764 15822
rect 1708 15148 1764 15204
rect 1708 14306 1764 14308
rect 1708 14254 1710 14306
rect 1710 14254 1762 14306
rect 1762 14254 1764 14306
rect 1708 14252 1764 14254
rect 1708 13468 1764 13524
rect 1708 11452 1764 11508
rect 1820 10780 1876 10836
rect 1708 10108 1764 10164
rect 2492 10780 2548 10836
rect 4732 16268 4788 16324
rect 3368 14922 3424 14924
rect 3368 14870 3370 14922
rect 3370 14870 3422 14922
rect 3422 14870 3424 14922
rect 3368 14868 3424 14870
rect 3472 14922 3528 14924
rect 3472 14870 3474 14922
rect 3474 14870 3526 14922
rect 3526 14870 3528 14922
rect 3472 14868 3528 14870
rect 3576 14922 3632 14924
rect 3576 14870 3578 14922
rect 3578 14870 3630 14922
rect 3630 14870 3632 14922
rect 3576 14868 3632 14870
rect 5964 16322 6020 16324
rect 5964 16270 5966 16322
rect 5966 16270 6018 16322
rect 6018 16270 6020 16322
rect 5964 16268 6020 16270
rect 5524 15706 5580 15708
rect 5524 15654 5526 15706
rect 5526 15654 5578 15706
rect 5578 15654 5580 15706
rect 5524 15652 5580 15654
rect 5628 15706 5684 15708
rect 5628 15654 5630 15706
rect 5630 15654 5682 15706
rect 5682 15654 5684 15706
rect 5628 15652 5684 15654
rect 5732 15706 5788 15708
rect 5732 15654 5734 15706
rect 5734 15654 5786 15706
rect 5786 15654 5788 15706
rect 5732 15652 5788 15654
rect 6636 16098 6692 16100
rect 6636 16046 6638 16098
rect 6638 16046 6690 16098
rect 6690 16046 6692 16098
rect 6636 16044 6692 16046
rect 7680 16490 7736 16492
rect 7680 16438 7682 16490
rect 7682 16438 7734 16490
rect 7734 16438 7736 16490
rect 7680 16436 7736 16438
rect 7784 16490 7840 16492
rect 7784 16438 7786 16490
rect 7786 16438 7838 16490
rect 7838 16438 7840 16490
rect 7784 16436 7840 16438
rect 7888 16490 7944 16492
rect 7888 16438 7890 16490
rect 7890 16438 7942 16490
rect 7942 16438 7944 16490
rect 7888 16436 7944 16438
rect 9100 16044 9156 16100
rect 7680 14922 7736 14924
rect 7680 14870 7682 14922
rect 7682 14870 7734 14922
rect 7734 14870 7736 14922
rect 7680 14868 7736 14870
rect 7784 14922 7840 14924
rect 7784 14870 7786 14922
rect 7786 14870 7838 14922
rect 7838 14870 7840 14922
rect 7784 14868 7840 14870
rect 7888 14922 7944 14924
rect 7888 14870 7890 14922
rect 7890 14870 7942 14922
rect 7942 14870 7944 14922
rect 7888 14868 7944 14870
rect 5524 14138 5580 14140
rect 5524 14086 5526 14138
rect 5526 14086 5578 14138
rect 5578 14086 5580 14138
rect 5524 14084 5580 14086
rect 5628 14138 5684 14140
rect 5628 14086 5630 14138
rect 5630 14086 5682 14138
rect 5682 14086 5684 14138
rect 5628 14084 5684 14086
rect 5732 14138 5788 14140
rect 5732 14086 5734 14138
rect 5734 14086 5786 14138
rect 5786 14086 5788 14138
rect 5732 14084 5788 14086
rect 4956 13468 5012 13524
rect 3368 13354 3424 13356
rect 3368 13302 3370 13354
rect 3370 13302 3422 13354
rect 3422 13302 3424 13354
rect 3368 13300 3424 13302
rect 3472 13354 3528 13356
rect 3472 13302 3474 13354
rect 3474 13302 3526 13354
rect 3526 13302 3528 13354
rect 3472 13300 3528 13302
rect 3576 13354 3632 13356
rect 3576 13302 3578 13354
rect 3578 13302 3630 13354
rect 3630 13302 3632 13354
rect 3576 13300 3632 13302
rect 5524 12570 5580 12572
rect 5524 12518 5526 12570
rect 5526 12518 5578 12570
rect 5578 12518 5580 12570
rect 5524 12516 5580 12518
rect 5628 12570 5684 12572
rect 5628 12518 5630 12570
rect 5630 12518 5682 12570
rect 5682 12518 5684 12570
rect 5628 12516 5684 12518
rect 5732 12570 5788 12572
rect 5732 12518 5734 12570
rect 5734 12518 5786 12570
rect 5786 12518 5788 12570
rect 5732 12516 5788 12518
rect 4956 12124 5012 12180
rect 3368 11786 3424 11788
rect 3368 11734 3370 11786
rect 3370 11734 3422 11786
rect 3422 11734 3424 11786
rect 3368 11732 3424 11734
rect 3472 11786 3528 11788
rect 3472 11734 3474 11786
rect 3474 11734 3526 11786
rect 3526 11734 3528 11786
rect 3472 11732 3528 11734
rect 3576 11786 3632 11788
rect 3576 11734 3578 11786
rect 3578 11734 3630 11786
rect 3630 11734 3632 11786
rect 3576 11732 3632 11734
rect 7680 13354 7736 13356
rect 7680 13302 7682 13354
rect 7682 13302 7734 13354
rect 7734 13302 7736 13354
rect 7680 13300 7736 13302
rect 7784 13354 7840 13356
rect 7784 13302 7786 13354
rect 7786 13302 7838 13354
rect 7838 13302 7840 13354
rect 7784 13300 7840 13302
rect 7888 13354 7944 13356
rect 7888 13302 7890 13354
rect 7890 13302 7942 13354
rect 7942 13302 7944 13354
rect 7888 13300 7944 13302
rect 8092 12236 8148 12292
rect 8988 13468 9044 13524
rect 6076 12012 6132 12068
rect 5180 11394 5236 11396
rect 5180 11342 5182 11394
rect 5182 11342 5234 11394
rect 5234 11342 5236 11394
rect 5180 11340 5236 11342
rect 5524 11002 5580 11004
rect 5524 10950 5526 11002
rect 5526 10950 5578 11002
rect 5578 10950 5580 11002
rect 5524 10948 5580 10950
rect 5628 11002 5684 11004
rect 5628 10950 5630 11002
rect 5630 10950 5682 11002
rect 5682 10950 5684 11002
rect 5628 10948 5684 10950
rect 5732 11002 5788 11004
rect 5732 10950 5734 11002
rect 5734 10950 5786 11002
rect 5786 10950 5788 11002
rect 5732 10948 5788 10950
rect 3368 10218 3424 10220
rect 3368 10166 3370 10218
rect 3370 10166 3422 10218
rect 3422 10166 3424 10218
rect 3368 10164 3424 10166
rect 3472 10218 3528 10220
rect 3472 10166 3474 10218
rect 3474 10166 3526 10218
rect 3526 10166 3528 10218
rect 3472 10164 3528 10166
rect 3576 10218 3632 10220
rect 3576 10166 3578 10218
rect 3578 10166 3630 10218
rect 3630 10166 3632 10218
rect 3576 10164 3632 10166
rect 3276 9996 3332 10052
rect 2044 9772 2100 9828
rect 6860 12066 6916 12068
rect 6860 12014 6862 12066
rect 6862 12014 6914 12066
rect 6914 12014 6916 12066
rect 6860 12012 6916 12014
rect 8316 11900 8372 11956
rect 7680 11786 7736 11788
rect 7680 11734 7682 11786
rect 7682 11734 7734 11786
rect 7734 11734 7736 11786
rect 7680 11732 7736 11734
rect 7784 11786 7840 11788
rect 7784 11734 7786 11786
rect 7786 11734 7838 11786
rect 7838 11734 7840 11786
rect 7784 11732 7840 11734
rect 7888 11786 7944 11788
rect 7888 11734 7890 11786
rect 7890 11734 7942 11786
rect 7942 11734 7944 11786
rect 7888 11732 7944 11734
rect 6412 11394 6468 11396
rect 6412 11342 6414 11394
rect 6414 11342 6466 11394
rect 6466 11342 6468 11394
rect 6412 11340 6468 11342
rect 8540 11116 8596 11172
rect 5516 9996 5572 10052
rect 9836 15706 9892 15708
rect 9836 15654 9838 15706
rect 9838 15654 9890 15706
rect 9890 15654 9892 15706
rect 9836 15652 9892 15654
rect 9940 15706 9996 15708
rect 9940 15654 9942 15706
rect 9942 15654 9994 15706
rect 9994 15654 9996 15706
rect 9940 15652 9996 15654
rect 10044 15706 10100 15708
rect 10044 15654 10046 15706
rect 10046 15654 10098 15706
rect 10098 15654 10100 15706
rect 10044 15652 10100 15654
rect 11992 16490 12048 16492
rect 11992 16438 11994 16490
rect 11994 16438 12046 16490
rect 12046 16438 12048 16490
rect 11992 16436 12048 16438
rect 12096 16490 12152 16492
rect 12096 16438 12098 16490
rect 12098 16438 12150 16490
rect 12150 16438 12152 16490
rect 12096 16436 12152 16438
rect 12200 16490 12256 16492
rect 12200 16438 12202 16490
rect 12202 16438 12254 16490
rect 12254 16438 12256 16490
rect 12200 16436 12256 16438
rect 16304 16490 16360 16492
rect 16304 16438 16306 16490
rect 16306 16438 16358 16490
rect 16358 16438 16360 16490
rect 16304 16436 16360 16438
rect 16408 16490 16464 16492
rect 16408 16438 16410 16490
rect 16410 16438 16462 16490
rect 16462 16438 16464 16490
rect 16408 16436 16464 16438
rect 16512 16490 16568 16492
rect 16512 16438 16514 16490
rect 16514 16438 16566 16490
rect 16566 16438 16568 16490
rect 16512 16436 16568 16438
rect 16156 15932 16212 15988
rect 16940 15986 16996 15988
rect 16940 15934 16942 15986
rect 16942 15934 16994 15986
rect 16994 15934 16996 15986
rect 16940 15932 16996 15934
rect 9836 14138 9892 14140
rect 9836 14086 9838 14138
rect 9838 14086 9890 14138
rect 9890 14086 9892 14138
rect 9836 14084 9892 14086
rect 9940 14138 9996 14140
rect 9940 14086 9942 14138
rect 9942 14086 9994 14138
rect 9994 14086 9996 14138
rect 9940 14084 9996 14086
rect 10044 14138 10100 14140
rect 10044 14086 10046 14138
rect 10046 14086 10098 14138
rect 10098 14086 10100 14138
rect 10044 14084 10100 14086
rect 9836 12570 9892 12572
rect 9836 12518 9838 12570
rect 9838 12518 9890 12570
rect 9890 12518 9892 12570
rect 9836 12516 9892 12518
rect 9940 12570 9996 12572
rect 9940 12518 9942 12570
rect 9942 12518 9994 12570
rect 9994 12518 9996 12570
rect 9940 12516 9996 12518
rect 10044 12570 10100 12572
rect 10044 12518 10046 12570
rect 10046 12518 10098 12570
rect 10098 12518 10100 12570
rect 10044 12516 10100 12518
rect 9884 12290 9940 12292
rect 9884 12238 9886 12290
rect 9886 12238 9938 12290
rect 9938 12238 9940 12290
rect 9884 12236 9940 12238
rect 10332 12290 10388 12292
rect 10332 12238 10334 12290
rect 10334 12238 10386 12290
rect 10386 12238 10388 12290
rect 10332 12236 10388 12238
rect 10220 11954 10276 11956
rect 10220 11902 10222 11954
rect 10222 11902 10274 11954
rect 10274 11902 10276 11954
rect 10220 11900 10276 11902
rect 9772 11116 9828 11172
rect 16380 15874 16436 15876
rect 16380 15822 16382 15874
rect 16382 15822 16434 15874
rect 16434 15822 16436 15874
rect 16380 15820 16436 15822
rect 14148 15706 14204 15708
rect 14148 15654 14150 15706
rect 14150 15654 14202 15706
rect 14202 15654 14204 15706
rect 14148 15652 14204 15654
rect 14252 15706 14308 15708
rect 14252 15654 14254 15706
rect 14254 15654 14306 15706
rect 14306 15654 14308 15706
rect 14252 15652 14308 15654
rect 14356 15706 14412 15708
rect 14356 15654 14358 15706
rect 14358 15654 14410 15706
rect 14410 15654 14412 15706
rect 14356 15652 14412 15654
rect 19516 15820 19572 15876
rect 18460 15706 18516 15708
rect 18460 15654 18462 15706
rect 18462 15654 18514 15706
rect 18514 15654 18516 15706
rect 18460 15652 18516 15654
rect 18564 15706 18620 15708
rect 18564 15654 18566 15706
rect 18566 15654 18618 15706
rect 18618 15654 18620 15706
rect 18564 15652 18620 15654
rect 18668 15706 18724 15708
rect 18668 15654 18670 15706
rect 18670 15654 18722 15706
rect 18722 15654 18724 15706
rect 18668 15652 18724 15654
rect 11992 14922 12048 14924
rect 11992 14870 11994 14922
rect 11994 14870 12046 14922
rect 12046 14870 12048 14922
rect 11992 14868 12048 14870
rect 12096 14922 12152 14924
rect 12096 14870 12098 14922
rect 12098 14870 12150 14922
rect 12150 14870 12152 14922
rect 12096 14868 12152 14870
rect 12200 14922 12256 14924
rect 12200 14870 12202 14922
rect 12202 14870 12254 14922
rect 12254 14870 12256 14922
rect 12200 14868 12256 14870
rect 16304 14922 16360 14924
rect 16304 14870 16306 14922
rect 16306 14870 16358 14922
rect 16358 14870 16360 14922
rect 16304 14868 16360 14870
rect 16408 14922 16464 14924
rect 16408 14870 16410 14922
rect 16410 14870 16462 14922
rect 16462 14870 16464 14922
rect 16408 14868 16464 14870
rect 16512 14922 16568 14924
rect 16512 14870 16514 14922
rect 16514 14870 16566 14922
rect 16566 14870 16568 14922
rect 16512 14868 16568 14870
rect 14148 14138 14204 14140
rect 14148 14086 14150 14138
rect 14150 14086 14202 14138
rect 14202 14086 14204 14138
rect 14148 14084 14204 14086
rect 14252 14138 14308 14140
rect 14252 14086 14254 14138
rect 14254 14086 14306 14138
rect 14306 14086 14308 14138
rect 14252 14084 14308 14086
rect 14356 14138 14412 14140
rect 14356 14086 14358 14138
rect 14358 14086 14410 14138
rect 14410 14086 14412 14138
rect 14356 14084 14412 14086
rect 18460 14138 18516 14140
rect 18460 14086 18462 14138
rect 18462 14086 18514 14138
rect 18514 14086 18516 14138
rect 18460 14084 18516 14086
rect 18564 14138 18620 14140
rect 18564 14086 18566 14138
rect 18566 14086 18618 14138
rect 18618 14086 18620 14138
rect 18564 14084 18620 14086
rect 18668 14138 18724 14140
rect 18668 14086 18670 14138
rect 18670 14086 18722 14138
rect 18722 14086 18724 14138
rect 18668 14084 18724 14086
rect 11992 13354 12048 13356
rect 11992 13302 11994 13354
rect 11994 13302 12046 13354
rect 12046 13302 12048 13354
rect 11992 13300 12048 13302
rect 12096 13354 12152 13356
rect 12096 13302 12098 13354
rect 12098 13302 12150 13354
rect 12150 13302 12152 13354
rect 12096 13300 12152 13302
rect 12200 13354 12256 13356
rect 12200 13302 12202 13354
rect 12202 13302 12254 13354
rect 12254 13302 12256 13354
rect 12200 13300 12256 13302
rect 16304 13354 16360 13356
rect 16304 13302 16306 13354
rect 16306 13302 16358 13354
rect 16358 13302 16360 13354
rect 16304 13300 16360 13302
rect 16408 13354 16464 13356
rect 16408 13302 16410 13354
rect 16410 13302 16462 13354
rect 16462 13302 16464 13354
rect 16408 13300 16464 13302
rect 16512 13354 16568 13356
rect 16512 13302 16514 13354
rect 16514 13302 16566 13354
rect 16566 13302 16568 13354
rect 16512 13300 16568 13302
rect 14148 12570 14204 12572
rect 14148 12518 14150 12570
rect 14150 12518 14202 12570
rect 14202 12518 14204 12570
rect 14148 12516 14204 12518
rect 14252 12570 14308 12572
rect 14252 12518 14254 12570
rect 14254 12518 14306 12570
rect 14306 12518 14308 12570
rect 14252 12516 14308 12518
rect 14356 12570 14412 12572
rect 14356 12518 14358 12570
rect 14358 12518 14410 12570
rect 14410 12518 14412 12570
rect 14356 12516 14412 12518
rect 18460 12570 18516 12572
rect 18460 12518 18462 12570
rect 18462 12518 18514 12570
rect 18514 12518 18516 12570
rect 18460 12516 18516 12518
rect 18564 12570 18620 12572
rect 18564 12518 18566 12570
rect 18566 12518 18618 12570
rect 18618 12518 18620 12570
rect 18564 12516 18620 12518
rect 18668 12570 18724 12572
rect 18668 12518 18670 12570
rect 18670 12518 18722 12570
rect 18722 12518 18724 12570
rect 18668 12516 18724 12518
rect 12236 12236 12292 12292
rect 11992 11786 12048 11788
rect 11992 11734 11994 11786
rect 11994 11734 12046 11786
rect 12046 11734 12048 11786
rect 11992 11732 12048 11734
rect 12096 11786 12152 11788
rect 12096 11734 12098 11786
rect 12098 11734 12150 11786
rect 12150 11734 12152 11786
rect 12096 11732 12152 11734
rect 12200 11786 12256 11788
rect 12200 11734 12202 11786
rect 12202 11734 12254 11786
rect 12254 11734 12256 11786
rect 12200 11732 12256 11734
rect 9836 11002 9892 11004
rect 9836 10950 9838 11002
rect 9838 10950 9890 11002
rect 9890 10950 9892 11002
rect 9836 10948 9892 10950
rect 9940 11002 9996 11004
rect 9940 10950 9942 11002
rect 9942 10950 9994 11002
rect 9994 10950 9996 11002
rect 9940 10948 9996 10950
rect 10044 11002 10100 11004
rect 10044 10950 10046 11002
rect 10046 10950 10098 11002
rect 10098 10950 10100 11002
rect 10044 10948 10100 10950
rect 7532 10444 7588 10500
rect 7680 10218 7736 10220
rect 7680 10166 7682 10218
rect 7682 10166 7734 10218
rect 7734 10166 7736 10218
rect 7680 10164 7736 10166
rect 7784 10218 7840 10220
rect 7784 10166 7786 10218
rect 7786 10166 7838 10218
rect 7838 10166 7840 10218
rect 7784 10164 7840 10166
rect 7888 10218 7944 10220
rect 7888 10166 7890 10218
rect 7890 10166 7942 10218
rect 7942 10166 7944 10218
rect 7888 10164 7944 10166
rect 6076 9548 6132 9604
rect 5524 9434 5580 9436
rect 5524 9382 5526 9434
rect 5526 9382 5578 9434
rect 5578 9382 5580 9434
rect 5524 9380 5580 9382
rect 5628 9434 5684 9436
rect 5628 9382 5630 9434
rect 5630 9382 5682 9434
rect 5682 9382 5684 9434
rect 5628 9380 5684 9382
rect 5732 9434 5788 9436
rect 5732 9382 5734 9434
rect 5734 9382 5786 9434
rect 5786 9382 5788 9434
rect 5732 9380 5788 9382
rect 3368 8650 3424 8652
rect 3368 8598 3370 8650
rect 3370 8598 3422 8650
rect 3422 8598 3424 8650
rect 3368 8596 3424 8598
rect 3472 8650 3528 8652
rect 3472 8598 3474 8650
rect 3474 8598 3526 8650
rect 3526 8598 3528 8650
rect 3472 8596 3528 8598
rect 3576 8650 3632 8652
rect 3576 8598 3578 8650
rect 3578 8598 3630 8650
rect 3630 8598 3632 8650
rect 3576 8596 3632 8598
rect 7420 9602 7476 9604
rect 7420 9550 7422 9602
rect 7422 9550 7474 9602
rect 7474 9550 7476 9602
rect 7420 9548 7476 9550
rect 7680 8650 7736 8652
rect 7680 8598 7682 8650
rect 7682 8598 7734 8650
rect 7734 8598 7736 8650
rect 7680 8596 7736 8598
rect 7784 8650 7840 8652
rect 7784 8598 7786 8650
rect 7786 8598 7838 8650
rect 7838 8598 7840 8650
rect 7784 8596 7840 8598
rect 7888 8650 7944 8652
rect 7888 8598 7890 8650
rect 7890 8598 7942 8650
rect 7942 8598 7944 8650
rect 7888 8596 7944 8598
rect 5628 8316 5684 8372
rect 6636 8370 6692 8372
rect 6636 8318 6638 8370
rect 6638 8318 6690 8370
rect 6690 8318 6692 8370
rect 6636 8316 6692 8318
rect 1708 8146 1764 8148
rect 1708 8094 1710 8146
rect 1710 8094 1762 8146
rect 1762 8094 1764 8146
rect 1708 8092 1764 8094
rect 2044 8034 2100 8036
rect 2044 7982 2046 8034
rect 2046 7982 2098 8034
rect 2098 7982 2100 8034
rect 2044 7980 2100 7982
rect 5524 7866 5580 7868
rect 5524 7814 5526 7866
rect 5526 7814 5578 7866
rect 5578 7814 5580 7866
rect 5524 7812 5580 7814
rect 5628 7866 5684 7868
rect 5628 7814 5630 7866
rect 5630 7814 5682 7866
rect 5682 7814 5684 7866
rect 5628 7812 5684 7814
rect 5732 7866 5788 7868
rect 5732 7814 5734 7866
rect 5734 7814 5786 7866
rect 5786 7814 5788 7866
rect 5732 7812 5788 7814
rect 2380 7420 2436 7476
rect 2828 7420 2884 7476
rect 1708 5404 1764 5460
rect 812 4956 868 5012
rect 28 3388 84 3444
rect 1708 4956 1764 5012
rect 2044 6412 2100 6468
rect 1932 5068 1988 5124
rect 2268 4956 2324 5012
rect 2380 4898 2436 4900
rect 2380 4846 2382 4898
rect 2382 4846 2434 4898
rect 2434 4846 2436 4898
rect 2380 4844 2436 4846
rect 2044 4562 2100 4564
rect 2044 4510 2046 4562
rect 2046 4510 2098 4562
rect 2098 4510 2100 4562
rect 2044 4508 2100 4510
rect 2268 4396 2324 4452
rect 3368 7082 3424 7084
rect 3368 7030 3370 7082
rect 3370 7030 3422 7082
rect 3422 7030 3424 7082
rect 3368 7028 3424 7030
rect 3472 7082 3528 7084
rect 3472 7030 3474 7082
rect 3474 7030 3526 7082
rect 3526 7030 3528 7082
rect 3472 7028 3528 7030
rect 3576 7082 3632 7084
rect 3576 7030 3578 7082
rect 3578 7030 3630 7082
rect 3630 7030 3632 7082
rect 3576 7028 3632 7030
rect 6748 6636 6804 6692
rect 2940 6524 2996 6580
rect 2380 3388 2436 3444
rect 5524 6298 5580 6300
rect 5524 6246 5526 6298
rect 5526 6246 5578 6298
rect 5578 6246 5580 6298
rect 5524 6244 5580 6246
rect 5628 6298 5684 6300
rect 5628 6246 5630 6298
rect 5630 6246 5682 6298
rect 5682 6246 5684 6298
rect 5628 6244 5684 6246
rect 5732 6298 5788 6300
rect 5732 6246 5734 6298
rect 5734 6246 5786 6298
rect 5786 6246 5788 6298
rect 5732 6244 5788 6246
rect 6076 5964 6132 6020
rect 3368 5514 3424 5516
rect 3368 5462 3370 5514
rect 3370 5462 3422 5514
rect 3422 5462 3424 5514
rect 3368 5460 3424 5462
rect 3472 5514 3528 5516
rect 3472 5462 3474 5514
rect 3474 5462 3526 5514
rect 3526 5462 3528 5514
rect 3472 5460 3528 5462
rect 3576 5514 3632 5516
rect 3576 5462 3578 5514
rect 3578 5462 3630 5514
rect 3630 5462 3632 5514
rect 3576 5460 3632 5462
rect 3612 5122 3668 5124
rect 3612 5070 3614 5122
rect 3614 5070 3666 5122
rect 3666 5070 3668 5122
rect 3612 5068 3668 5070
rect 4956 4956 5012 5012
rect 3052 4060 3108 4116
rect 3368 3946 3424 3948
rect 3368 3894 3370 3946
rect 3370 3894 3422 3946
rect 3422 3894 3424 3946
rect 3368 3892 3424 3894
rect 3472 3946 3528 3948
rect 3472 3894 3474 3946
rect 3474 3894 3526 3946
rect 3526 3894 3528 3946
rect 3472 3892 3528 3894
rect 3576 3946 3632 3948
rect 3576 3894 3578 3946
rect 3578 3894 3630 3946
rect 3630 3894 3632 3946
rect 3576 3892 3632 3894
rect 3612 3388 3668 3444
rect 4284 3948 4340 4004
rect 5964 4844 6020 4900
rect 5524 4730 5580 4732
rect 5524 4678 5526 4730
rect 5526 4678 5578 4730
rect 5578 4678 5580 4730
rect 5524 4676 5580 4678
rect 5628 4730 5684 4732
rect 5628 4678 5630 4730
rect 5630 4678 5682 4730
rect 5682 4678 5684 4730
rect 5628 4676 5684 4678
rect 5732 4730 5788 4732
rect 5732 4678 5734 4730
rect 5734 4678 5786 4730
rect 5786 4678 5788 4730
rect 5732 4676 5788 4678
rect 5524 3162 5580 3164
rect 5524 3110 5526 3162
rect 5526 3110 5578 3162
rect 5578 3110 5580 3162
rect 5524 3108 5580 3110
rect 5628 3162 5684 3164
rect 5628 3110 5630 3162
rect 5630 3110 5682 3162
rect 5682 3110 5684 3162
rect 5628 3108 5684 3110
rect 5732 3162 5788 3164
rect 5732 3110 5734 3162
rect 5734 3110 5786 3162
rect 5786 3110 5788 3162
rect 5732 3108 5788 3110
rect 7084 6018 7140 6020
rect 7084 5966 7086 6018
rect 7086 5966 7138 6018
rect 7138 5966 7140 6018
rect 7084 5964 7140 5966
rect 7420 6412 7476 6468
rect 7680 7082 7736 7084
rect 7680 7030 7682 7082
rect 7682 7030 7734 7082
rect 7734 7030 7736 7082
rect 7680 7028 7736 7030
rect 7784 7082 7840 7084
rect 7784 7030 7786 7082
rect 7786 7030 7838 7082
rect 7838 7030 7840 7082
rect 7784 7028 7840 7030
rect 7888 7082 7944 7084
rect 7888 7030 7890 7082
rect 7890 7030 7942 7082
rect 7942 7030 7944 7082
rect 7888 7028 7944 7030
rect 9100 9884 9156 9940
rect 9100 9266 9156 9268
rect 9100 9214 9102 9266
rect 9102 9214 9154 9266
rect 9154 9214 9156 9266
rect 9100 9212 9156 9214
rect 9660 9996 9716 10052
rect 9996 10386 10052 10388
rect 9996 10334 9998 10386
rect 9998 10334 10050 10386
rect 10050 10334 10052 10386
rect 9996 10332 10052 10334
rect 9884 9548 9940 9604
rect 10332 10220 10388 10276
rect 9836 9434 9892 9436
rect 9836 9382 9838 9434
rect 9838 9382 9890 9434
rect 9890 9382 9892 9434
rect 9836 9380 9892 9382
rect 9940 9434 9996 9436
rect 9940 9382 9942 9434
rect 9942 9382 9994 9434
rect 9994 9382 9996 9434
rect 9940 9380 9996 9382
rect 10044 9434 10100 9436
rect 10044 9382 10046 9434
rect 10046 9382 10098 9434
rect 10098 9382 10100 9434
rect 10044 9380 10100 9382
rect 9836 7866 9892 7868
rect 9836 7814 9838 7866
rect 9838 7814 9890 7866
rect 9890 7814 9892 7866
rect 9836 7812 9892 7814
rect 9940 7866 9996 7868
rect 9940 7814 9942 7866
rect 9942 7814 9994 7866
rect 9994 7814 9996 7866
rect 9940 7812 9996 7814
rect 10044 7866 10100 7868
rect 10044 7814 10046 7866
rect 10046 7814 10098 7866
rect 10098 7814 10100 7866
rect 10044 7812 10100 7814
rect 10892 10498 10948 10500
rect 10892 10446 10894 10498
rect 10894 10446 10946 10498
rect 10946 10446 10948 10498
rect 10892 10444 10948 10446
rect 10556 10332 10612 10388
rect 10556 9212 10612 9268
rect 8428 7474 8484 7476
rect 8428 7422 8430 7474
rect 8430 7422 8482 7474
rect 8482 7422 8484 7474
rect 8428 7420 8484 7422
rect 8204 6690 8260 6692
rect 8204 6638 8206 6690
rect 8206 6638 8258 6690
rect 8258 6638 8260 6690
rect 8204 6636 8260 6638
rect 8092 5906 8148 5908
rect 8092 5854 8094 5906
rect 8094 5854 8146 5906
rect 8146 5854 8148 5906
rect 8092 5852 8148 5854
rect 7680 5514 7736 5516
rect 7680 5462 7682 5514
rect 7682 5462 7734 5514
rect 7734 5462 7736 5514
rect 7680 5460 7736 5462
rect 7784 5514 7840 5516
rect 7784 5462 7786 5514
rect 7786 5462 7838 5514
rect 7838 5462 7840 5514
rect 7784 5460 7840 5462
rect 7888 5514 7944 5516
rect 7888 5462 7890 5514
rect 7890 5462 7942 5514
rect 7942 5462 7944 5514
rect 7888 5460 7944 5462
rect 7308 4508 7364 4564
rect 8092 4620 8148 4676
rect 7680 3946 7736 3948
rect 7680 3894 7682 3946
rect 7682 3894 7734 3946
rect 7734 3894 7736 3946
rect 7680 3892 7736 3894
rect 7784 3946 7840 3948
rect 7784 3894 7786 3946
rect 7786 3894 7838 3946
rect 7838 3894 7840 3946
rect 7784 3892 7840 3894
rect 7888 3946 7944 3948
rect 7888 3894 7890 3946
rect 7890 3894 7942 3946
rect 7942 3894 7944 3946
rect 7888 3892 7944 3894
rect 8316 5794 8372 5796
rect 8316 5742 8318 5794
rect 8318 5742 8370 5794
rect 8370 5742 8372 5794
rect 8316 5740 8372 5742
rect 8428 5068 8484 5124
rect 8540 5852 8596 5908
rect 8428 4620 8484 4676
rect 8652 4956 8708 5012
rect 8540 4396 8596 4452
rect 8988 5404 9044 5460
rect 9100 4226 9156 4228
rect 9100 4174 9102 4226
rect 9102 4174 9154 4226
rect 9154 4174 9156 4226
rect 9100 4172 9156 4174
rect 9996 6636 10052 6692
rect 9548 5122 9604 5124
rect 9548 5070 9550 5122
rect 9550 5070 9602 5122
rect 9602 5070 9604 5122
rect 9548 5068 9604 5070
rect 9836 6298 9892 6300
rect 9836 6246 9838 6298
rect 9838 6246 9890 6298
rect 9890 6246 9892 6298
rect 9836 6244 9892 6246
rect 9940 6298 9996 6300
rect 9940 6246 9942 6298
rect 9942 6246 9994 6298
rect 9994 6246 9996 6298
rect 9940 6244 9996 6246
rect 10044 6298 10100 6300
rect 10044 6246 10046 6298
rect 10046 6246 10098 6298
rect 10098 6246 10100 6298
rect 10044 6244 10100 6246
rect 10220 6188 10276 6244
rect 9836 4730 9892 4732
rect 9836 4678 9838 4730
rect 9838 4678 9890 4730
rect 9890 4678 9892 4730
rect 9836 4676 9892 4678
rect 9940 4730 9996 4732
rect 9940 4678 9942 4730
rect 9942 4678 9994 4730
rect 9994 4678 9996 4730
rect 9940 4676 9996 4678
rect 10044 4730 10100 4732
rect 10044 4678 10046 4730
rect 10046 4678 10098 4730
rect 10098 4678 10100 4730
rect 10044 4676 10100 4678
rect 10332 5740 10388 5796
rect 10444 5682 10500 5684
rect 10444 5630 10446 5682
rect 10446 5630 10498 5682
rect 10498 5630 10500 5682
rect 10444 5628 10500 5630
rect 10444 5404 10500 5460
rect 10220 4396 10276 4452
rect 9436 3724 9492 3780
rect 9884 4172 9940 4228
rect 11992 10218 12048 10220
rect 11992 10166 11994 10218
rect 11994 10166 12046 10218
rect 12046 10166 12048 10218
rect 11992 10164 12048 10166
rect 12096 10218 12152 10220
rect 12096 10166 12098 10218
rect 12098 10166 12150 10218
rect 12150 10166 12152 10218
rect 12096 10164 12152 10166
rect 12200 10218 12256 10220
rect 12200 10166 12202 10218
rect 12202 10166 12254 10218
rect 12254 10166 12256 10218
rect 12200 10164 12256 10166
rect 11676 9996 11732 10052
rect 16304 11786 16360 11788
rect 16304 11734 16306 11786
rect 16306 11734 16358 11786
rect 16358 11734 16360 11786
rect 16304 11732 16360 11734
rect 16408 11786 16464 11788
rect 16408 11734 16410 11786
rect 16410 11734 16462 11786
rect 16462 11734 16464 11786
rect 16408 11732 16464 11734
rect 16512 11786 16568 11788
rect 16512 11734 16514 11786
rect 16514 11734 16566 11786
rect 16566 11734 16568 11786
rect 16512 11732 16568 11734
rect 14148 11002 14204 11004
rect 14148 10950 14150 11002
rect 14150 10950 14202 11002
rect 14202 10950 14204 11002
rect 14148 10948 14204 10950
rect 14252 11002 14308 11004
rect 14252 10950 14254 11002
rect 14254 10950 14306 11002
rect 14306 10950 14308 11002
rect 14252 10948 14308 10950
rect 14356 11002 14412 11004
rect 14356 10950 14358 11002
rect 14358 10950 14410 11002
rect 14410 10950 14412 11002
rect 14356 10948 14412 10950
rect 18460 11002 18516 11004
rect 18460 10950 18462 11002
rect 18462 10950 18514 11002
rect 18514 10950 18516 11002
rect 18460 10948 18516 10950
rect 18564 11002 18620 11004
rect 18564 10950 18566 11002
rect 18566 10950 18618 11002
rect 18618 10950 18620 11002
rect 18564 10948 18620 10950
rect 18668 11002 18724 11004
rect 18668 10950 18670 11002
rect 18670 10950 18722 11002
rect 18722 10950 18724 11002
rect 18668 10948 18724 10950
rect 12572 10386 12628 10388
rect 12572 10334 12574 10386
rect 12574 10334 12626 10386
rect 12626 10334 12628 10386
rect 12572 10332 12628 10334
rect 11228 9212 11284 9268
rect 16304 10218 16360 10220
rect 16304 10166 16306 10218
rect 16306 10166 16358 10218
rect 16358 10166 16360 10218
rect 16304 10164 16360 10166
rect 16408 10218 16464 10220
rect 16408 10166 16410 10218
rect 16410 10166 16462 10218
rect 16462 10166 16464 10218
rect 16408 10164 16464 10166
rect 16512 10218 16568 10220
rect 16512 10166 16514 10218
rect 16514 10166 16566 10218
rect 16566 10166 16568 10218
rect 16512 10164 16568 10166
rect 13468 9996 13524 10052
rect 12796 9772 12852 9828
rect 10780 6578 10836 6580
rect 10780 6526 10782 6578
rect 10782 6526 10834 6578
rect 10834 6526 10836 6578
rect 10780 6524 10836 6526
rect 10556 4172 10612 4228
rect 10668 6076 10724 6132
rect 9884 3276 9940 3332
rect 9436 3164 9492 3220
rect 9836 3162 9892 3164
rect 9836 3110 9838 3162
rect 9838 3110 9890 3162
rect 9890 3110 9892 3162
rect 9836 3108 9892 3110
rect 9940 3162 9996 3164
rect 9940 3110 9942 3162
rect 9942 3110 9994 3162
rect 9994 3110 9996 3162
rect 9940 3108 9996 3110
rect 10044 3162 10100 3164
rect 10044 3110 10046 3162
rect 10046 3110 10098 3162
rect 10098 3110 10100 3162
rect 10044 3108 10100 3110
rect 10668 3388 10724 3444
rect 10892 4060 10948 4116
rect 13692 9772 13748 9828
rect 12460 9714 12516 9716
rect 12460 9662 12462 9714
rect 12462 9662 12514 9714
rect 12514 9662 12516 9714
rect 12460 9660 12516 9662
rect 13580 9714 13636 9716
rect 13580 9662 13582 9714
rect 13582 9662 13634 9714
rect 13634 9662 13636 9714
rect 13580 9660 13636 9662
rect 11788 9548 11844 9604
rect 12684 9100 12740 9156
rect 11564 4844 11620 4900
rect 11452 3500 11508 3556
rect 11992 8650 12048 8652
rect 11992 8598 11994 8650
rect 11994 8598 12046 8650
rect 12046 8598 12048 8650
rect 11992 8596 12048 8598
rect 12096 8650 12152 8652
rect 12096 8598 12098 8650
rect 12098 8598 12150 8650
rect 12150 8598 12152 8650
rect 12096 8596 12152 8598
rect 12200 8650 12256 8652
rect 12200 8598 12202 8650
rect 12202 8598 12254 8650
rect 12254 8598 12256 8650
rect 12200 8596 12256 8598
rect 11992 7082 12048 7084
rect 11992 7030 11994 7082
rect 11994 7030 12046 7082
rect 12046 7030 12048 7082
rect 11992 7028 12048 7030
rect 12096 7082 12152 7084
rect 12096 7030 12098 7082
rect 12098 7030 12150 7082
rect 12150 7030 12152 7082
rect 12096 7028 12152 7030
rect 12200 7082 12256 7084
rect 12200 7030 12202 7082
rect 12202 7030 12254 7082
rect 12254 7030 12256 7082
rect 12200 7028 12256 7030
rect 12012 6018 12068 6020
rect 12012 5966 12014 6018
rect 12014 5966 12066 6018
rect 12066 5966 12068 6018
rect 12012 5964 12068 5966
rect 11992 5514 12048 5516
rect 11992 5462 11994 5514
rect 11994 5462 12046 5514
rect 12046 5462 12048 5514
rect 11992 5460 12048 5462
rect 12096 5514 12152 5516
rect 12096 5462 12098 5514
rect 12098 5462 12150 5514
rect 12150 5462 12152 5514
rect 12096 5460 12152 5462
rect 12200 5514 12256 5516
rect 12200 5462 12202 5514
rect 12202 5462 12254 5514
rect 12254 5462 12256 5514
rect 12200 5460 12256 5462
rect 12684 7980 12740 8036
rect 12572 6690 12628 6692
rect 12572 6638 12574 6690
rect 12574 6638 12626 6690
rect 12626 6638 12628 6690
rect 12572 6636 12628 6638
rect 13468 9154 13524 9156
rect 13468 9102 13470 9154
rect 13470 9102 13522 9154
rect 13522 9102 13524 9154
rect 13468 9100 13524 9102
rect 12572 5906 12628 5908
rect 12572 5854 12574 5906
rect 12574 5854 12626 5906
rect 12626 5854 12628 5906
rect 12572 5852 12628 5854
rect 12460 5516 12516 5572
rect 12460 4956 12516 5012
rect 11992 3946 12048 3948
rect 11992 3894 11994 3946
rect 11994 3894 12046 3946
rect 12046 3894 12048 3946
rect 11992 3892 12048 3894
rect 12096 3946 12152 3948
rect 12096 3894 12098 3946
rect 12098 3894 12150 3946
rect 12150 3894 12152 3946
rect 12096 3892 12152 3894
rect 12200 3946 12256 3948
rect 12200 3894 12202 3946
rect 12202 3894 12254 3946
rect 12254 3894 12256 3946
rect 12200 3892 12256 3894
rect 11900 3554 11956 3556
rect 11900 3502 11902 3554
rect 11902 3502 11954 3554
rect 11954 3502 11956 3554
rect 11900 3500 11956 3502
rect 12684 3554 12740 3556
rect 12684 3502 12686 3554
rect 12686 3502 12738 3554
rect 12738 3502 12740 3554
rect 12684 3500 12740 3502
rect 12796 3388 12852 3444
rect 14148 9434 14204 9436
rect 14148 9382 14150 9434
rect 14150 9382 14202 9434
rect 14202 9382 14204 9434
rect 14148 9380 14204 9382
rect 14252 9434 14308 9436
rect 14252 9382 14254 9434
rect 14254 9382 14306 9434
rect 14306 9382 14308 9434
rect 14252 9380 14308 9382
rect 14356 9434 14412 9436
rect 14356 9382 14358 9434
rect 14358 9382 14410 9434
rect 14410 9382 14412 9434
rect 14356 9380 14412 9382
rect 18460 9434 18516 9436
rect 18460 9382 18462 9434
rect 18462 9382 18514 9434
rect 18514 9382 18516 9434
rect 18460 9380 18516 9382
rect 18564 9434 18620 9436
rect 18564 9382 18566 9434
rect 18566 9382 18618 9434
rect 18618 9382 18620 9434
rect 18564 9380 18620 9382
rect 18668 9434 18724 9436
rect 18668 9382 18670 9434
rect 18670 9382 18722 9434
rect 18722 9382 18724 9434
rect 18668 9380 18724 9382
rect 13916 8204 13972 8260
rect 14148 7866 14204 7868
rect 14148 7814 14150 7866
rect 14150 7814 14202 7866
rect 14202 7814 14204 7866
rect 14148 7812 14204 7814
rect 14252 7866 14308 7868
rect 14252 7814 14254 7866
rect 14254 7814 14306 7866
rect 14306 7814 14308 7866
rect 14252 7812 14308 7814
rect 14356 7866 14412 7868
rect 14356 7814 14358 7866
rect 14358 7814 14410 7866
rect 14410 7814 14412 7866
rect 14356 7812 14412 7814
rect 17612 8764 17668 8820
rect 16304 8650 16360 8652
rect 16304 8598 16306 8650
rect 16306 8598 16358 8650
rect 16358 8598 16360 8650
rect 16304 8596 16360 8598
rect 16408 8650 16464 8652
rect 16408 8598 16410 8650
rect 16410 8598 16462 8650
rect 16462 8598 16464 8650
rect 16408 8596 16464 8598
rect 16512 8650 16568 8652
rect 16512 8598 16514 8650
rect 16514 8598 16566 8650
rect 16566 8598 16568 8650
rect 16512 8596 16568 8598
rect 18172 8764 18228 8820
rect 14700 8092 14756 8148
rect 17164 8204 17220 8260
rect 17836 8146 17892 8148
rect 17836 8094 17838 8146
rect 17838 8094 17890 8146
rect 17890 8094 17892 8146
rect 17836 8092 17892 8094
rect 17724 7474 17780 7476
rect 17724 7422 17726 7474
rect 17726 7422 17778 7474
rect 17778 7422 17780 7474
rect 17724 7420 17780 7422
rect 16304 7082 16360 7084
rect 16304 7030 16306 7082
rect 16306 7030 16358 7082
rect 16358 7030 16360 7082
rect 16304 7028 16360 7030
rect 16408 7082 16464 7084
rect 16408 7030 16410 7082
rect 16410 7030 16462 7082
rect 16462 7030 16464 7082
rect 16408 7028 16464 7030
rect 16512 7082 16568 7084
rect 16512 7030 16514 7082
rect 16514 7030 16566 7082
rect 16566 7030 16568 7082
rect 16512 7028 16568 7030
rect 14148 6298 14204 6300
rect 14148 6246 14150 6298
rect 14150 6246 14202 6298
rect 14202 6246 14204 6298
rect 14148 6244 14204 6246
rect 14252 6298 14308 6300
rect 14252 6246 14254 6298
rect 14254 6246 14306 6298
rect 14306 6246 14308 6298
rect 14252 6244 14308 6246
rect 14356 6298 14412 6300
rect 14356 6246 14358 6298
rect 14358 6246 14410 6298
rect 14410 6246 14412 6298
rect 14356 6244 14412 6246
rect 13356 3554 13412 3556
rect 13356 3502 13358 3554
rect 13358 3502 13410 3554
rect 13410 3502 13412 3554
rect 13356 3500 13412 3502
rect 13580 3388 13636 3444
rect 14148 4730 14204 4732
rect 14148 4678 14150 4730
rect 14150 4678 14202 4730
rect 14202 4678 14204 4730
rect 14148 4676 14204 4678
rect 14252 4730 14308 4732
rect 14252 4678 14254 4730
rect 14254 4678 14306 4730
rect 14306 4678 14308 4730
rect 14252 4676 14308 4678
rect 14356 4730 14412 4732
rect 14356 4678 14358 4730
rect 14358 4678 14410 4730
rect 14410 4678 14412 4730
rect 14356 4676 14412 4678
rect 14140 3442 14196 3444
rect 14140 3390 14142 3442
rect 14142 3390 14194 3442
rect 14194 3390 14196 3442
rect 14140 3388 14196 3390
rect 18172 8146 18228 8148
rect 18172 8094 18174 8146
rect 18174 8094 18226 8146
rect 18226 8094 18228 8146
rect 18172 8092 18228 8094
rect 18460 7866 18516 7868
rect 18460 7814 18462 7866
rect 18462 7814 18514 7866
rect 18514 7814 18516 7866
rect 18460 7812 18516 7814
rect 18564 7866 18620 7868
rect 18564 7814 18566 7866
rect 18566 7814 18618 7866
rect 18618 7814 18620 7866
rect 18564 7812 18620 7814
rect 18668 7866 18724 7868
rect 18668 7814 18670 7866
rect 18670 7814 18722 7866
rect 18722 7814 18724 7866
rect 18668 7812 18724 7814
rect 18460 6298 18516 6300
rect 18460 6246 18462 6298
rect 18462 6246 18514 6298
rect 18514 6246 18516 6298
rect 18460 6244 18516 6246
rect 18564 6298 18620 6300
rect 18564 6246 18566 6298
rect 18566 6246 18618 6298
rect 18618 6246 18620 6298
rect 18564 6244 18620 6246
rect 18668 6298 18724 6300
rect 18668 6246 18670 6298
rect 18670 6246 18722 6298
rect 18722 6246 18724 6298
rect 18668 6244 18724 6246
rect 17948 5964 18004 6020
rect 14588 4508 14644 4564
rect 15148 5852 15204 5908
rect 14148 3162 14204 3164
rect 14148 3110 14150 3162
rect 14150 3110 14202 3162
rect 14202 3110 14204 3162
rect 14148 3108 14204 3110
rect 14252 3162 14308 3164
rect 14252 3110 14254 3162
rect 14254 3110 14306 3162
rect 14306 3110 14308 3162
rect 14252 3108 14308 3110
rect 14356 3162 14412 3164
rect 14356 3110 14358 3162
rect 14358 3110 14410 3162
rect 14410 3110 14412 3162
rect 14356 3108 14412 3110
rect 14812 3500 14868 3556
rect 14924 3388 14980 3444
rect 16044 5516 16100 5572
rect 15708 4562 15764 4564
rect 15708 4510 15710 4562
rect 15710 4510 15762 4562
rect 15762 4510 15764 4562
rect 15708 4508 15764 4510
rect 15484 3554 15540 3556
rect 15484 3502 15486 3554
rect 15486 3502 15538 3554
rect 15538 3502 15540 3554
rect 15484 3500 15540 3502
rect 15372 3388 15428 3444
rect 16304 5514 16360 5516
rect 16304 5462 16306 5514
rect 16306 5462 16358 5514
rect 16358 5462 16360 5514
rect 16304 5460 16360 5462
rect 16408 5514 16464 5516
rect 16408 5462 16410 5514
rect 16410 5462 16462 5514
rect 16462 5462 16464 5514
rect 16408 5460 16464 5462
rect 16512 5514 16568 5516
rect 16512 5462 16514 5514
rect 16514 5462 16566 5514
rect 16566 5462 16568 5514
rect 16512 5460 16568 5462
rect 16492 4956 16548 5012
rect 16304 3946 16360 3948
rect 16304 3894 16306 3946
rect 16306 3894 16358 3946
rect 16358 3894 16360 3946
rect 16304 3892 16360 3894
rect 16408 3946 16464 3948
rect 16408 3894 16410 3946
rect 16410 3894 16462 3946
rect 16462 3894 16464 3946
rect 16408 3892 16464 3894
rect 16512 3946 16568 3948
rect 16512 3894 16514 3946
rect 16514 3894 16566 3946
rect 16566 3894 16568 3946
rect 16512 3892 16568 3894
rect 16044 3388 16100 3444
rect 16268 3388 16324 3444
rect 16828 4338 16884 4340
rect 16828 4286 16830 4338
rect 16830 4286 16882 4338
rect 16882 4286 16884 4338
rect 16828 4284 16884 4286
rect 17164 4284 17220 4340
rect 16716 3388 16772 3444
rect 16940 3724 16996 3780
rect 17164 3388 17220 3444
rect 17836 5628 17892 5684
rect 17724 4450 17780 4452
rect 17724 4398 17726 4450
rect 17726 4398 17778 4450
rect 17778 4398 17780 4450
rect 17724 4396 17780 4398
rect 17612 4172 17668 4228
rect 18060 4284 18116 4340
rect 18460 4730 18516 4732
rect 18460 4678 18462 4730
rect 18462 4678 18514 4730
rect 18514 4678 18516 4730
rect 18460 4676 18516 4678
rect 18564 4730 18620 4732
rect 18564 4678 18566 4730
rect 18566 4678 18618 4730
rect 18618 4678 18620 4730
rect 18564 4676 18620 4678
rect 18668 4730 18724 4732
rect 18668 4678 18670 4730
rect 18670 4678 18722 4730
rect 18722 4678 18724 4730
rect 18668 4676 18724 4678
rect 18460 3162 18516 3164
rect 18460 3110 18462 3162
rect 18462 3110 18514 3162
rect 18514 3110 18516 3162
rect 18460 3108 18516 3110
rect 18564 3162 18620 3164
rect 18564 3110 18566 3162
rect 18566 3110 18618 3162
rect 18618 3110 18620 3162
rect 18564 3108 18620 3110
rect 18668 3162 18724 3164
rect 18668 3110 18670 3162
rect 18670 3110 18722 3162
rect 18722 3110 18724 3162
rect 18668 3108 18724 3110
<< metal3 >>
rect 0 19488 800 19600
rect 19200 19488 20000 19600
rect 0 18816 800 18928
rect 19200 18816 20000 18928
rect 0 18144 800 18256
rect 19200 18144 20000 18256
rect 0 17472 800 17584
rect 19200 17472 20000 17584
rect 19200 16800 20000 16912
rect 3358 16436 3368 16492
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3632 16436 3642 16492
rect 7670 16436 7680 16492
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7944 16436 7954 16492
rect 11982 16436 11992 16492
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 12256 16436 12266 16492
rect 16294 16436 16304 16492
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16568 16436 16578 16492
rect 4722 16268 4732 16324
rect 4788 16268 5964 16324
rect 6020 16268 6030 16324
rect 19200 16128 20000 16240
rect 6626 16044 6636 16100
rect 6692 16044 9100 16100
rect 9156 16044 9166 16100
rect 16146 15932 16156 15988
rect 16212 15932 16940 15988
rect 16996 15932 17006 15988
rect 1698 15820 1708 15876
rect 1764 15820 1774 15876
rect 16370 15820 16380 15876
rect 16436 15820 19516 15876
rect 19572 15820 19582 15876
rect 0 15540 800 15568
rect 1708 15540 1764 15820
rect 5514 15652 5524 15708
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5788 15652 5798 15708
rect 9826 15652 9836 15708
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 10100 15652 10110 15708
rect 14138 15652 14148 15708
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14412 15652 14422 15708
rect 18450 15652 18460 15708
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18724 15652 18734 15708
rect 0 15484 1764 15540
rect 0 15456 800 15484
rect 19200 15456 20000 15568
rect 1698 15148 1708 15204
rect 1764 15148 1774 15204
rect 0 14868 800 14896
rect 1708 14868 1764 15148
rect 3358 14868 3368 14924
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3632 14868 3642 14924
rect 7670 14868 7680 14924
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7944 14868 7954 14924
rect 11982 14868 11992 14924
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 12256 14868 12266 14924
rect 16294 14868 16304 14924
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16568 14868 16578 14924
rect 0 14812 1764 14868
rect 0 14784 800 14812
rect 19200 14784 20000 14896
rect 1698 14252 1708 14308
rect 1764 14252 1774 14308
rect 0 14196 800 14224
rect 1708 14196 1764 14252
rect 0 14140 1764 14196
rect 0 14112 800 14140
rect 5514 14084 5524 14140
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5788 14084 5798 14140
rect 9826 14084 9836 14140
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 10100 14084 10110 14140
rect 14138 14084 14148 14140
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14412 14084 14422 14140
rect 18450 14084 18460 14140
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18724 14084 18734 14140
rect 19200 14112 20000 14224
rect 0 13524 800 13552
rect 0 13468 1708 13524
rect 1764 13468 1774 13524
rect 4946 13468 4956 13524
rect 5012 13468 8988 13524
rect 9044 13468 9054 13524
rect 0 13440 800 13468
rect 19200 13440 20000 13552
rect 3358 13300 3368 13356
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3632 13300 3642 13356
rect 7670 13300 7680 13356
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7944 13300 7954 13356
rect 11982 13300 11992 13356
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 12256 13300 12266 13356
rect 16294 13300 16304 13356
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16568 13300 16578 13356
rect 19200 12768 20000 12880
rect 5514 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5798 12572
rect 9826 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10110 12572
rect 14138 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14422 12572
rect 18450 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18734 12572
rect 8082 12236 8092 12292
rect 8148 12236 9884 12292
rect 9940 12236 10332 12292
rect 10388 12236 12236 12292
rect 12292 12236 12302 12292
rect 0 12180 800 12208
rect 0 12124 4956 12180
rect 5012 12124 5022 12180
rect 0 12096 800 12124
rect 19200 12096 20000 12208
rect 6066 12012 6076 12068
rect 6132 12012 6860 12068
rect 6916 12012 6926 12068
rect 8306 11900 8316 11956
rect 8372 11900 10220 11956
rect 10276 11900 10286 11956
rect 3358 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3642 11788
rect 7670 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7954 11788
rect 11982 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12266 11788
rect 16294 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16578 11788
rect 0 11508 800 11536
rect 0 11452 1708 11508
rect 1764 11452 1774 11508
rect 0 11424 800 11452
rect 19200 11424 20000 11536
rect 5170 11340 5180 11396
rect 5236 11340 6412 11396
rect 6468 11340 6478 11396
rect 8530 11116 8540 11172
rect 8596 11116 9772 11172
rect 9828 11116 9838 11172
rect 5514 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5798 11004
rect 9826 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10110 11004
rect 14138 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14422 11004
rect 18450 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18734 11004
rect 0 10836 800 10864
rect 0 10780 1820 10836
rect 1876 10780 2492 10836
rect 2548 10780 2558 10836
rect 0 10752 800 10780
rect 19200 10752 20000 10864
rect 7522 10444 7532 10500
rect 7588 10444 10892 10500
rect 10948 10444 10958 10500
rect 9986 10332 9996 10388
rect 10052 10332 10556 10388
rect 10612 10332 10622 10388
rect 11116 10332 12572 10388
rect 12628 10332 12638 10388
rect 11116 10276 11172 10332
rect 10322 10220 10332 10276
rect 10388 10220 11172 10276
rect 0 10164 800 10192
rect 3358 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3642 10220
rect 7670 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7954 10220
rect 11982 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12266 10220
rect 16294 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16578 10220
rect 0 10108 1708 10164
rect 1764 10108 1774 10164
rect 0 10080 800 10108
rect 19200 10080 20000 10192
rect 3266 9996 3276 10052
rect 3332 9940 3388 10052
rect 5506 9996 5516 10052
rect 5572 9996 9660 10052
rect 9716 9996 9726 10052
rect 11666 9996 11676 10052
rect 11732 9996 13468 10052
rect 13524 9996 13534 10052
rect 3332 9884 9100 9940
rect 9156 9884 9166 9940
rect 2034 9772 2044 9828
rect 2100 9772 3388 9828
rect 12786 9772 12796 9828
rect 12852 9772 13692 9828
rect 13748 9772 13758 9828
rect 3332 9716 3388 9772
rect 3332 9660 12460 9716
rect 12516 9660 13580 9716
rect 13636 9660 13646 9716
rect 6066 9548 6076 9604
rect 6132 9548 7420 9604
rect 7476 9548 7486 9604
rect 9874 9548 9884 9604
rect 9940 9548 11788 9604
rect 11844 9548 11854 9604
rect 5514 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5798 9436
rect 9826 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10110 9436
rect 14138 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14422 9436
rect 18450 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18734 9436
rect 19200 9408 20000 9520
rect 9090 9212 9100 9268
rect 9156 9212 10556 9268
rect 10612 9212 11228 9268
rect 11284 9212 11294 9268
rect 12674 9100 12684 9156
rect 12740 9100 13468 9156
rect 13524 9100 13534 9156
rect 19200 8820 20000 8848
rect 17602 8764 17612 8820
rect 17668 8764 18172 8820
rect 18228 8764 20000 8820
rect 19200 8736 20000 8764
rect 3358 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3642 8652
rect 7670 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7954 8652
rect 11982 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12266 8652
rect 16294 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16578 8652
rect 5618 8316 5628 8372
rect 5684 8316 6636 8372
rect 6692 8316 6702 8372
rect 13906 8204 13916 8260
rect 13972 8204 17164 8260
rect 17220 8204 17230 8260
rect 0 8148 800 8176
rect 19200 8148 20000 8176
rect 0 8092 1708 8148
rect 1764 8092 1774 8148
rect 14690 8092 14700 8148
rect 14756 8092 17836 8148
rect 17892 8092 17902 8148
rect 18162 8092 18172 8148
rect 18228 8092 20000 8148
rect 0 8064 800 8092
rect 19200 8064 20000 8092
rect 2034 7980 2044 8036
rect 2100 7980 12684 8036
rect 12740 7980 12750 8036
rect 5514 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5798 7868
rect 9826 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10110 7868
rect 14138 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14422 7868
rect 18450 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18734 7868
rect 0 7476 800 7504
rect 19200 7476 20000 7504
rect 0 7420 2380 7476
rect 2436 7420 2446 7476
rect 2818 7420 2828 7476
rect 2884 7420 8428 7476
rect 8484 7420 8494 7476
rect 17714 7420 17724 7476
rect 17780 7420 20000 7476
rect 0 7392 800 7420
rect 19200 7392 20000 7420
rect 3358 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3642 7084
rect 7670 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7954 7084
rect 11982 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12266 7084
rect 16294 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16578 7084
rect 19200 6720 20000 6832
rect 6738 6636 6748 6692
rect 6804 6636 8204 6692
rect 8260 6636 8270 6692
rect 9986 6636 9996 6692
rect 10052 6636 12572 6692
rect 12628 6636 12638 6692
rect 2930 6524 2940 6580
rect 2996 6524 10780 6580
rect 10836 6524 10846 6580
rect 2034 6412 2044 6468
rect 2100 6412 7420 6468
rect 7476 6412 7486 6468
rect 5514 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5798 6300
rect 9826 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10110 6300
rect 14138 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14422 6300
rect 18450 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18734 6300
rect 10210 6188 10220 6244
rect 10276 6188 10724 6244
rect 10668 6132 10724 6188
rect 10658 6076 10668 6132
rect 10724 6076 10734 6132
rect 19200 6048 20000 6160
rect 6066 5964 6076 6020
rect 6132 5964 7084 6020
rect 7140 5964 7150 6020
rect 12002 5964 12012 6020
rect 12068 5964 17948 6020
rect 18004 5964 18014 6020
rect 8082 5852 8092 5908
rect 8148 5852 8540 5908
rect 8596 5852 8606 5908
rect 12562 5852 12572 5908
rect 12628 5852 15148 5908
rect 15204 5852 15214 5908
rect 8306 5740 8316 5796
rect 8372 5740 10332 5796
rect 10388 5740 10398 5796
rect 10434 5628 10444 5684
rect 10500 5628 17836 5684
rect 17892 5628 17902 5684
rect 12450 5516 12460 5572
rect 12516 5516 16044 5572
rect 16100 5516 16110 5572
rect 0 5460 800 5488
rect 3358 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3642 5516
rect 7670 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7954 5516
rect 11982 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12266 5516
rect 16294 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16578 5516
rect 0 5404 1708 5460
rect 1764 5404 1774 5460
rect 8978 5404 8988 5460
rect 9044 5404 10444 5460
rect 10500 5404 10510 5460
rect 0 5376 800 5404
rect 19200 5376 20000 5488
rect 1922 5068 1932 5124
rect 1988 5068 3612 5124
rect 3668 5068 3678 5124
rect 8418 5068 8428 5124
rect 8484 5068 9548 5124
rect 9604 5068 9614 5124
rect 802 4956 812 5012
rect 868 4956 1708 5012
rect 1764 4956 2268 5012
rect 2324 4956 2334 5012
rect 4946 4956 4956 5012
rect 5012 4956 8652 5012
rect 8708 4956 8718 5012
rect 12450 4956 12460 5012
rect 12516 4956 16492 5012
rect 16548 4956 16558 5012
rect 2370 4844 2380 4900
rect 2436 4844 2446 4900
rect 5954 4844 5964 4900
rect 6020 4844 11564 4900
rect 11620 4844 11630 4900
rect 0 4788 800 4816
rect 2380 4788 2436 4844
rect 0 4732 2436 4788
rect 0 4704 800 4732
rect 5514 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5798 4732
rect 9826 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10110 4732
rect 14138 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14422 4732
rect 18450 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18734 4732
rect 19200 4704 20000 4816
rect 8082 4620 8092 4676
rect 8148 4620 8428 4676
rect 8484 4620 8494 4676
rect 2034 4508 2044 4564
rect 2100 4508 7308 4564
rect 7364 4508 7374 4564
rect 14578 4508 14588 4564
rect 14644 4508 15708 4564
rect 15764 4508 15774 4564
rect 2258 4396 2268 4452
rect 2324 4396 8540 4452
rect 8596 4396 8606 4452
rect 10210 4396 10220 4452
rect 10276 4396 17724 4452
rect 17780 4396 17790 4452
rect 16818 4284 16828 4340
rect 16884 4284 17164 4340
rect 17220 4284 18060 4340
rect 18116 4284 18126 4340
rect 9090 4172 9100 4228
rect 9156 4172 9884 4228
rect 9940 4172 9950 4228
rect 10546 4172 10556 4228
rect 10612 4172 17612 4228
rect 17668 4172 17678 4228
rect 0 4116 800 4144
rect 0 4060 3052 4116
rect 3108 4060 3118 4116
rect 4284 4060 10892 4116
rect 10948 4060 10958 4116
rect 0 4032 800 4060
rect 4284 4004 4340 4060
rect 19200 4032 20000 4144
rect 4274 3948 4284 4004
rect 4340 3948 4350 4004
rect 3358 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3642 3948
rect 7670 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7954 3948
rect 11982 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12266 3948
rect 16294 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16578 3948
rect 9426 3724 9436 3780
rect 9492 3724 16940 3780
rect 16996 3724 17006 3780
rect 11442 3500 11452 3556
rect 11508 3500 11900 3556
rect 11956 3500 11966 3556
rect 12674 3500 12684 3556
rect 12740 3500 13356 3556
rect 13412 3500 13422 3556
rect 14802 3500 14812 3556
rect 14868 3500 15484 3556
rect 15540 3500 15550 3556
rect 18 3388 28 3444
rect 84 3388 2380 3444
rect 2436 3388 2446 3444
rect 3602 3388 3612 3444
rect 3668 3388 10668 3444
rect 10724 3388 10734 3444
rect 12786 3388 12796 3444
rect 12852 3388 13580 3444
rect 13636 3388 14140 3444
rect 14196 3388 14206 3444
rect 14914 3388 14924 3444
rect 14980 3388 15372 3444
rect 15428 3388 16044 3444
rect 16100 3388 16110 3444
rect 16258 3388 16268 3444
rect 16324 3388 16716 3444
rect 16772 3388 17164 3444
rect 17220 3388 17230 3444
rect 19200 3360 20000 3472
rect 9436 3276 9884 3332
rect 9940 3276 9950 3332
rect 9436 3220 9492 3276
rect 9426 3164 9436 3220
rect 9492 3164 9502 3220
rect 5514 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5798 3164
rect 9826 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10110 3164
rect 14138 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14422 3164
rect 18450 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18734 3164
rect 19200 2688 20000 2800
rect 19200 2016 20000 2128
rect 19200 1344 20000 1456
rect 19200 672 20000 784
rect 19200 0 20000 112
<< via3 >>
rect 3368 16436 3424 16492
rect 3472 16436 3528 16492
rect 3576 16436 3632 16492
rect 7680 16436 7736 16492
rect 7784 16436 7840 16492
rect 7888 16436 7944 16492
rect 11992 16436 12048 16492
rect 12096 16436 12152 16492
rect 12200 16436 12256 16492
rect 16304 16436 16360 16492
rect 16408 16436 16464 16492
rect 16512 16436 16568 16492
rect 5524 15652 5580 15708
rect 5628 15652 5684 15708
rect 5732 15652 5788 15708
rect 9836 15652 9892 15708
rect 9940 15652 9996 15708
rect 10044 15652 10100 15708
rect 14148 15652 14204 15708
rect 14252 15652 14308 15708
rect 14356 15652 14412 15708
rect 18460 15652 18516 15708
rect 18564 15652 18620 15708
rect 18668 15652 18724 15708
rect 3368 14868 3424 14924
rect 3472 14868 3528 14924
rect 3576 14868 3632 14924
rect 7680 14868 7736 14924
rect 7784 14868 7840 14924
rect 7888 14868 7944 14924
rect 11992 14868 12048 14924
rect 12096 14868 12152 14924
rect 12200 14868 12256 14924
rect 16304 14868 16360 14924
rect 16408 14868 16464 14924
rect 16512 14868 16568 14924
rect 5524 14084 5580 14140
rect 5628 14084 5684 14140
rect 5732 14084 5788 14140
rect 9836 14084 9892 14140
rect 9940 14084 9996 14140
rect 10044 14084 10100 14140
rect 14148 14084 14204 14140
rect 14252 14084 14308 14140
rect 14356 14084 14412 14140
rect 18460 14084 18516 14140
rect 18564 14084 18620 14140
rect 18668 14084 18724 14140
rect 3368 13300 3424 13356
rect 3472 13300 3528 13356
rect 3576 13300 3632 13356
rect 7680 13300 7736 13356
rect 7784 13300 7840 13356
rect 7888 13300 7944 13356
rect 11992 13300 12048 13356
rect 12096 13300 12152 13356
rect 12200 13300 12256 13356
rect 16304 13300 16360 13356
rect 16408 13300 16464 13356
rect 16512 13300 16568 13356
rect 5524 12516 5580 12572
rect 5628 12516 5684 12572
rect 5732 12516 5788 12572
rect 9836 12516 9892 12572
rect 9940 12516 9996 12572
rect 10044 12516 10100 12572
rect 14148 12516 14204 12572
rect 14252 12516 14308 12572
rect 14356 12516 14412 12572
rect 18460 12516 18516 12572
rect 18564 12516 18620 12572
rect 18668 12516 18724 12572
rect 3368 11732 3424 11788
rect 3472 11732 3528 11788
rect 3576 11732 3632 11788
rect 7680 11732 7736 11788
rect 7784 11732 7840 11788
rect 7888 11732 7944 11788
rect 11992 11732 12048 11788
rect 12096 11732 12152 11788
rect 12200 11732 12256 11788
rect 16304 11732 16360 11788
rect 16408 11732 16464 11788
rect 16512 11732 16568 11788
rect 5524 10948 5580 11004
rect 5628 10948 5684 11004
rect 5732 10948 5788 11004
rect 9836 10948 9892 11004
rect 9940 10948 9996 11004
rect 10044 10948 10100 11004
rect 14148 10948 14204 11004
rect 14252 10948 14308 11004
rect 14356 10948 14412 11004
rect 18460 10948 18516 11004
rect 18564 10948 18620 11004
rect 18668 10948 18724 11004
rect 3368 10164 3424 10220
rect 3472 10164 3528 10220
rect 3576 10164 3632 10220
rect 7680 10164 7736 10220
rect 7784 10164 7840 10220
rect 7888 10164 7944 10220
rect 11992 10164 12048 10220
rect 12096 10164 12152 10220
rect 12200 10164 12256 10220
rect 16304 10164 16360 10220
rect 16408 10164 16464 10220
rect 16512 10164 16568 10220
rect 5524 9380 5580 9436
rect 5628 9380 5684 9436
rect 5732 9380 5788 9436
rect 9836 9380 9892 9436
rect 9940 9380 9996 9436
rect 10044 9380 10100 9436
rect 14148 9380 14204 9436
rect 14252 9380 14308 9436
rect 14356 9380 14412 9436
rect 18460 9380 18516 9436
rect 18564 9380 18620 9436
rect 18668 9380 18724 9436
rect 3368 8596 3424 8652
rect 3472 8596 3528 8652
rect 3576 8596 3632 8652
rect 7680 8596 7736 8652
rect 7784 8596 7840 8652
rect 7888 8596 7944 8652
rect 11992 8596 12048 8652
rect 12096 8596 12152 8652
rect 12200 8596 12256 8652
rect 16304 8596 16360 8652
rect 16408 8596 16464 8652
rect 16512 8596 16568 8652
rect 5524 7812 5580 7868
rect 5628 7812 5684 7868
rect 5732 7812 5788 7868
rect 9836 7812 9892 7868
rect 9940 7812 9996 7868
rect 10044 7812 10100 7868
rect 14148 7812 14204 7868
rect 14252 7812 14308 7868
rect 14356 7812 14412 7868
rect 18460 7812 18516 7868
rect 18564 7812 18620 7868
rect 18668 7812 18724 7868
rect 3368 7028 3424 7084
rect 3472 7028 3528 7084
rect 3576 7028 3632 7084
rect 7680 7028 7736 7084
rect 7784 7028 7840 7084
rect 7888 7028 7944 7084
rect 11992 7028 12048 7084
rect 12096 7028 12152 7084
rect 12200 7028 12256 7084
rect 16304 7028 16360 7084
rect 16408 7028 16464 7084
rect 16512 7028 16568 7084
rect 5524 6244 5580 6300
rect 5628 6244 5684 6300
rect 5732 6244 5788 6300
rect 9836 6244 9892 6300
rect 9940 6244 9996 6300
rect 10044 6244 10100 6300
rect 14148 6244 14204 6300
rect 14252 6244 14308 6300
rect 14356 6244 14412 6300
rect 18460 6244 18516 6300
rect 18564 6244 18620 6300
rect 18668 6244 18724 6300
rect 3368 5460 3424 5516
rect 3472 5460 3528 5516
rect 3576 5460 3632 5516
rect 7680 5460 7736 5516
rect 7784 5460 7840 5516
rect 7888 5460 7944 5516
rect 11992 5460 12048 5516
rect 12096 5460 12152 5516
rect 12200 5460 12256 5516
rect 16304 5460 16360 5516
rect 16408 5460 16464 5516
rect 16512 5460 16568 5516
rect 5524 4676 5580 4732
rect 5628 4676 5684 4732
rect 5732 4676 5788 4732
rect 9836 4676 9892 4732
rect 9940 4676 9996 4732
rect 10044 4676 10100 4732
rect 14148 4676 14204 4732
rect 14252 4676 14308 4732
rect 14356 4676 14412 4732
rect 18460 4676 18516 4732
rect 18564 4676 18620 4732
rect 18668 4676 18724 4732
rect 3368 3892 3424 3948
rect 3472 3892 3528 3948
rect 3576 3892 3632 3948
rect 7680 3892 7736 3948
rect 7784 3892 7840 3948
rect 7888 3892 7944 3948
rect 11992 3892 12048 3948
rect 12096 3892 12152 3948
rect 12200 3892 12256 3948
rect 16304 3892 16360 3948
rect 16408 3892 16464 3948
rect 16512 3892 16568 3948
rect 5524 3108 5580 3164
rect 5628 3108 5684 3164
rect 5732 3108 5788 3164
rect 9836 3108 9892 3164
rect 9940 3108 9996 3164
rect 10044 3108 10100 3164
rect 14148 3108 14204 3164
rect 14252 3108 14308 3164
rect 14356 3108 14412 3164
rect 18460 3108 18516 3164
rect 18564 3108 18620 3164
rect 18668 3108 18724 3164
<< metal4 >>
rect 3340 16492 3660 16524
rect 3340 16436 3368 16492
rect 3424 16436 3472 16492
rect 3528 16436 3576 16492
rect 3632 16436 3660 16492
rect 3340 14924 3660 16436
rect 3340 14868 3368 14924
rect 3424 14868 3472 14924
rect 3528 14868 3576 14924
rect 3632 14868 3660 14924
rect 3340 13356 3660 14868
rect 3340 13300 3368 13356
rect 3424 13300 3472 13356
rect 3528 13300 3576 13356
rect 3632 13300 3660 13356
rect 3340 11788 3660 13300
rect 3340 11732 3368 11788
rect 3424 11732 3472 11788
rect 3528 11732 3576 11788
rect 3632 11732 3660 11788
rect 3340 10220 3660 11732
rect 3340 10164 3368 10220
rect 3424 10164 3472 10220
rect 3528 10164 3576 10220
rect 3632 10164 3660 10220
rect 3340 8652 3660 10164
rect 3340 8596 3368 8652
rect 3424 8596 3472 8652
rect 3528 8596 3576 8652
rect 3632 8596 3660 8652
rect 3340 7084 3660 8596
rect 3340 7028 3368 7084
rect 3424 7028 3472 7084
rect 3528 7028 3576 7084
rect 3632 7028 3660 7084
rect 3340 5516 3660 7028
rect 3340 5460 3368 5516
rect 3424 5460 3472 5516
rect 3528 5460 3576 5516
rect 3632 5460 3660 5516
rect 3340 3948 3660 5460
rect 3340 3892 3368 3948
rect 3424 3892 3472 3948
rect 3528 3892 3576 3948
rect 3632 3892 3660 3948
rect 3340 3076 3660 3892
rect 5496 15708 5816 16524
rect 5496 15652 5524 15708
rect 5580 15652 5628 15708
rect 5684 15652 5732 15708
rect 5788 15652 5816 15708
rect 5496 14140 5816 15652
rect 5496 14084 5524 14140
rect 5580 14084 5628 14140
rect 5684 14084 5732 14140
rect 5788 14084 5816 14140
rect 5496 12572 5816 14084
rect 5496 12516 5524 12572
rect 5580 12516 5628 12572
rect 5684 12516 5732 12572
rect 5788 12516 5816 12572
rect 5496 11004 5816 12516
rect 5496 10948 5524 11004
rect 5580 10948 5628 11004
rect 5684 10948 5732 11004
rect 5788 10948 5816 11004
rect 5496 9436 5816 10948
rect 5496 9380 5524 9436
rect 5580 9380 5628 9436
rect 5684 9380 5732 9436
rect 5788 9380 5816 9436
rect 5496 7868 5816 9380
rect 5496 7812 5524 7868
rect 5580 7812 5628 7868
rect 5684 7812 5732 7868
rect 5788 7812 5816 7868
rect 5496 6300 5816 7812
rect 5496 6244 5524 6300
rect 5580 6244 5628 6300
rect 5684 6244 5732 6300
rect 5788 6244 5816 6300
rect 5496 4732 5816 6244
rect 5496 4676 5524 4732
rect 5580 4676 5628 4732
rect 5684 4676 5732 4732
rect 5788 4676 5816 4732
rect 5496 3164 5816 4676
rect 5496 3108 5524 3164
rect 5580 3108 5628 3164
rect 5684 3108 5732 3164
rect 5788 3108 5816 3164
rect 5496 3076 5816 3108
rect 7652 16492 7972 16524
rect 7652 16436 7680 16492
rect 7736 16436 7784 16492
rect 7840 16436 7888 16492
rect 7944 16436 7972 16492
rect 7652 14924 7972 16436
rect 7652 14868 7680 14924
rect 7736 14868 7784 14924
rect 7840 14868 7888 14924
rect 7944 14868 7972 14924
rect 7652 13356 7972 14868
rect 7652 13300 7680 13356
rect 7736 13300 7784 13356
rect 7840 13300 7888 13356
rect 7944 13300 7972 13356
rect 7652 11788 7972 13300
rect 7652 11732 7680 11788
rect 7736 11732 7784 11788
rect 7840 11732 7888 11788
rect 7944 11732 7972 11788
rect 7652 10220 7972 11732
rect 7652 10164 7680 10220
rect 7736 10164 7784 10220
rect 7840 10164 7888 10220
rect 7944 10164 7972 10220
rect 7652 8652 7972 10164
rect 7652 8596 7680 8652
rect 7736 8596 7784 8652
rect 7840 8596 7888 8652
rect 7944 8596 7972 8652
rect 7652 7084 7972 8596
rect 7652 7028 7680 7084
rect 7736 7028 7784 7084
rect 7840 7028 7888 7084
rect 7944 7028 7972 7084
rect 7652 5516 7972 7028
rect 7652 5460 7680 5516
rect 7736 5460 7784 5516
rect 7840 5460 7888 5516
rect 7944 5460 7972 5516
rect 7652 3948 7972 5460
rect 7652 3892 7680 3948
rect 7736 3892 7784 3948
rect 7840 3892 7888 3948
rect 7944 3892 7972 3948
rect 7652 3076 7972 3892
rect 9808 15708 10128 16524
rect 9808 15652 9836 15708
rect 9892 15652 9940 15708
rect 9996 15652 10044 15708
rect 10100 15652 10128 15708
rect 9808 14140 10128 15652
rect 9808 14084 9836 14140
rect 9892 14084 9940 14140
rect 9996 14084 10044 14140
rect 10100 14084 10128 14140
rect 9808 12572 10128 14084
rect 9808 12516 9836 12572
rect 9892 12516 9940 12572
rect 9996 12516 10044 12572
rect 10100 12516 10128 12572
rect 9808 11004 10128 12516
rect 9808 10948 9836 11004
rect 9892 10948 9940 11004
rect 9996 10948 10044 11004
rect 10100 10948 10128 11004
rect 9808 9436 10128 10948
rect 9808 9380 9836 9436
rect 9892 9380 9940 9436
rect 9996 9380 10044 9436
rect 10100 9380 10128 9436
rect 9808 7868 10128 9380
rect 9808 7812 9836 7868
rect 9892 7812 9940 7868
rect 9996 7812 10044 7868
rect 10100 7812 10128 7868
rect 9808 6300 10128 7812
rect 9808 6244 9836 6300
rect 9892 6244 9940 6300
rect 9996 6244 10044 6300
rect 10100 6244 10128 6300
rect 9808 4732 10128 6244
rect 9808 4676 9836 4732
rect 9892 4676 9940 4732
rect 9996 4676 10044 4732
rect 10100 4676 10128 4732
rect 9808 3164 10128 4676
rect 9808 3108 9836 3164
rect 9892 3108 9940 3164
rect 9996 3108 10044 3164
rect 10100 3108 10128 3164
rect 9808 3076 10128 3108
rect 11964 16492 12284 16524
rect 11964 16436 11992 16492
rect 12048 16436 12096 16492
rect 12152 16436 12200 16492
rect 12256 16436 12284 16492
rect 11964 14924 12284 16436
rect 11964 14868 11992 14924
rect 12048 14868 12096 14924
rect 12152 14868 12200 14924
rect 12256 14868 12284 14924
rect 11964 13356 12284 14868
rect 11964 13300 11992 13356
rect 12048 13300 12096 13356
rect 12152 13300 12200 13356
rect 12256 13300 12284 13356
rect 11964 11788 12284 13300
rect 11964 11732 11992 11788
rect 12048 11732 12096 11788
rect 12152 11732 12200 11788
rect 12256 11732 12284 11788
rect 11964 10220 12284 11732
rect 11964 10164 11992 10220
rect 12048 10164 12096 10220
rect 12152 10164 12200 10220
rect 12256 10164 12284 10220
rect 11964 8652 12284 10164
rect 11964 8596 11992 8652
rect 12048 8596 12096 8652
rect 12152 8596 12200 8652
rect 12256 8596 12284 8652
rect 11964 7084 12284 8596
rect 11964 7028 11992 7084
rect 12048 7028 12096 7084
rect 12152 7028 12200 7084
rect 12256 7028 12284 7084
rect 11964 5516 12284 7028
rect 11964 5460 11992 5516
rect 12048 5460 12096 5516
rect 12152 5460 12200 5516
rect 12256 5460 12284 5516
rect 11964 3948 12284 5460
rect 11964 3892 11992 3948
rect 12048 3892 12096 3948
rect 12152 3892 12200 3948
rect 12256 3892 12284 3948
rect 11964 3076 12284 3892
rect 14120 15708 14440 16524
rect 14120 15652 14148 15708
rect 14204 15652 14252 15708
rect 14308 15652 14356 15708
rect 14412 15652 14440 15708
rect 14120 14140 14440 15652
rect 14120 14084 14148 14140
rect 14204 14084 14252 14140
rect 14308 14084 14356 14140
rect 14412 14084 14440 14140
rect 14120 12572 14440 14084
rect 14120 12516 14148 12572
rect 14204 12516 14252 12572
rect 14308 12516 14356 12572
rect 14412 12516 14440 12572
rect 14120 11004 14440 12516
rect 14120 10948 14148 11004
rect 14204 10948 14252 11004
rect 14308 10948 14356 11004
rect 14412 10948 14440 11004
rect 14120 9436 14440 10948
rect 14120 9380 14148 9436
rect 14204 9380 14252 9436
rect 14308 9380 14356 9436
rect 14412 9380 14440 9436
rect 14120 7868 14440 9380
rect 14120 7812 14148 7868
rect 14204 7812 14252 7868
rect 14308 7812 14356 7868
rect 14412 7812 14440 7868
rect 14120 6300 14440 7812
rect 14120 6244 14148 6300
rect 14204 6244 14252 6300
rect 14308 6244 14356 6300
rect 14412 6244 14440 6300
rect 14120 4732 14440 6244
rect 14120 4676 14148 4732
rect 14204 4676 14252 4732
rect 14308 4676 14356 4732
rect 14412 4676 14440 4732
rect 14120 3164 14440 4676
rect 14120 3108 14148 3164
rect 14204 3108 14252 3164
rect 14308 3108 14356 3164
rect 14412 3108 14440 3164
rect 14120 3076 14440 3108
rect 16276 16492 16596 16524
rect 16276 16436 16304 16492
rect 16360 16436 16408 16492
rect 16464 16436 16512 16492
rect 16568 16436 16596 16492
rect 16276 14924 16596 16436
rect 16276 14868 16304 14924
rect 16360 14868 16408 14924
rect 16464 14868 16512 14924
rect 16568 14868 16596 14924
rect 16276 13356 16596 14868
rect 16276 13300 16304 13356
rect 16360 13300 16408 13356
rect 16464 13300 16512 13356
rect 16568 13300 16596 13356
rect 16276 11788 16596 13300
rect 16276 11732 16304 11788
rect 16360 11732 16408 11788
rect 16464 11732 16512 11788
rect 16568 11732 16596 11788
rect 16276 10220 16596 11732
rect 16276 10164 16304 10220
rect 16360 10164 16408 10220
rect 16464 10164 16512 10220
rect 16568 10164 16596 10220
rect 16276 8652 16596 10164
rect 16276 8596 16304 8652
rect 16360 8596 16408 8652
rect 16464 8596 16512 8652
rect 16568 8596 16596 8652
rect 16276 7084 16596 8596
rect 16276 7028 16304 7084
rect 16360 7028 16408 7084
rect 16464 7028 16512 7084
rect 16568 7028 16596 7084
rect 16276 5516 16596 7028
rect 16276 5460 16304 5516
rect 16360 5460 16408 5516
rect 16464 5460 16512 5516
rect 16568 5460 16596 5516
rect 16276 3948 16596 5460
rect 16276 3892 16304 3948
rect 16360 3892 16408 3948
rect 16464 3892 16512 3948
rect 16568 3892 16596 3948
rect 16276 3076 16596 3892
rect 18432 15708 18752 16524
rect 18432 15652 18460 15708
rect 18516 15652 18564 15708
rect 18620 15652 18668 15708
rect 18724 15652 18752 15708
rect 18432 14140 18752 15652
rect 18432 14084 18460 14140
rect 18516 14084 18564 14140
rect 18620 14084 18668 14140
rect 18724 14084 18752 14140
rect 18432 12572 18752 14084
rect 18432 12516 18460 12572
rect 18516 12516 18564 12572
rect 18620 12516 18668 12572
rect 18724 12516 18752 12572
rect 18432 11004 18752 12516
rect 18432 10948 18460 11004
rect 18516 10948 18564 11004
rect 18620 10948 18668 11004
rect 18724 10948 18752 11004
rect 18432 9436 18752 10948
rect 18432 9380 18460 9436
rect 18516 9380 18564 9436
rect 18620 9380 18668 9436
rect 18724 9380 18752 9436
rect 18432 7868 18752 9380
rect 18432 7812 18460 7868
rect 18516 7812 18564 7868
rect 18620 7812 18668 7868
rect 18724 7812 18752 7868
rect 18432 6300 18752 7812
rect 18432 6244 18460 6300
rect 18516 6244 18564 6300
rect 18620 6244 18668 6300
rect 18724 6244 18752 6300
rect 18432 4732 18752 6244
rect 18432 4676 18460 4732
rect 18516 4676 18564 4732
rect 18620 4676 18668 4732
rect 18724 4676 18752 4732
rect 18432 3164 18752 4676
rect 18432 3108 18460 3164
rect 18516 3108 18564 3164
rect 18620 3108 18668 3164
rect 18724 3108 18752 3164
rect 18432 3076 18752 3108
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _24_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10416 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _25_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _26_
timestamp 1698431365
transform -1 0 13104 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _27_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14784 0 -1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _28_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 14896 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _29_
timestamp 1698431365
transform -1 0 10640 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _30_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11088 0 -1 9408
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _31_
timestamp 1698431365
transform 1 0 9744 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _32_
timestamp 1698431365
transform 1 0 7168 0 -1 7840
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _33_
timestamp 1698431365
transform 1 0 6944 0 -1 6272
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _34_
timestamp 1698431365
transform 1 0 8064 0 1 6272
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _35_
timestamp 1698431365
transform 1 0 7952 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _36_
timestamp 1698431365
transform 1 0 9408 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _37_
timestamp 1698431365
transform 1 0 10416 0 -1 7840
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _38_
timestamp 1698431365
transform -1 0 13888 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _39_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 10640 0 -1 10976
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _40_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 7952 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _41_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 10080 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _42_
timestamp 1698431365
transform -1 0 10528 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _43_
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _44_
timestamp 1698431365
transform 1 0 12320 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _45_
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _46_
timestamp 1698431365
transform 1 0 5600 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _47_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 -1 9408
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  _48__71 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__dffrnq_1  _48_
timestamp 1698431365
transform 1 0 5376 0 -1 10976
box -86 -86 3894 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _49_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5936 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 7504 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 18368 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform 1 0 2688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 10192 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform 1 0 2240 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform 1 0 1792 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform 1 0 3808 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform 1 0 3136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform 1 0 4816 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform 1 0 6944 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 5488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 4368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 17696 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform 1 0 8064 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform 1 0 7616 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 15008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input17_I
timestamp 1698431365
transform -1 0 17696 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input18_I
timestamp 1698431365
transform -1 0 14336 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input19_I
timestamp 1698431365
transform -1 0 15568 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input20_I
timestamp 1698431365
transform -1 0 13664 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input21_I
timestamp 1698431365
transform -1 0 15680 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input22_I
timestamp 1698431365
transform 1 0 17696 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input23_I
timestamp 1698431365
transform -1 0 18368 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input24_I
timestamp 1698431365
transform -1 0 17248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input25_I
timestamp 1698431365
transform -1 0 17696 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input26_I
timestamp 1698431365
transform -1 0 16800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input27_I
timestamp 1698431365
transform -1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input28_I
timestamp 1698431365
transform -1 0 10864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input29_I
timestamp 1698431365
transform -1 0 11536 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input30_I
timestamp 1698431365
transform 1 0 3584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input31_I
timestamp 1698431365
transform -1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input32_I
timestamp 1698431365
transform 1 0 6384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input33_I
timestamp 1698431365
transform -1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input34_I
timestamp 1698431365
transform -1 0 10864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input35_I
timestamp 1698431365
transform 1 0 1792 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input36_I
timestamp 1698431365
transform 1 0 2464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 6272 0 1 10976
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_wb_clk_i
timestamp 1698431365
transform -1 0 11872 0 1 7840
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_wb_clk_i
timestamp 1698431365
transform -1 0 11312 0 1 14112
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_36
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_70
timestamp 1698431365
transform 1 0 9184 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_72 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 9408 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_97
timestamp 1698431365
transform 1 0 12208 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_99
timestamp 1698431365
transform 1 0 12432 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_134
timestamp 1698431365
transform 1 0 16352 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_150
timestamp 1698431365
transform 1 0 18144 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_18 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_24
timestamp 1698431365
transform 1 0 4032 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_26
timestamp 1698431365
transform 1 0 4256 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_29
timestamp 1698431365
transform 1 0 4592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_33
timestamp 1698431365
transform 1 0 5040 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_43
timestamp 1698431365
transform 1 0 6160 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_47
timestamp 1698431365
transform 1 0 6608 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_49
timestamp 1698431365
transform 1 0 6832 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_52
timestamp 1698431365
transform 1 0 7168 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_58
timestamp 1698431365
transform 1 0 7840 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_62
timestamp 1698431365
transform 1 0 8288 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_66
timestamp 1698431365
transform 1 0 8736 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_76
timestamp 1698431365
transform 1 0 9856 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_79
timestamp 1698431365
transform 1 0 10192 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_85
timestamp 1698431365
transform 1 0 10864 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_91 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 11536 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_107
timestamp 1698431365
transform 1 0 13328 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_110
timestamp 1698431365
transform 1 0 13664 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_116
timestamp 1698431365
transform 1 0 14336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_122
timestamp 1698431365
transform 1 0 15008 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_124
timestamp 1698431365
transform 1 0 15232 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_133
timestamp 1698431365
transform 1 0 16240 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698431365
transform 1 0 17472 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_151
timestamp 1698431365
transform 1 0 18256 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_12
timestamp 1698431365
transform 1 0 2688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_18
timestamp 1698431365
transform 1 0 3360 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_22 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_30
timestamp 1698431365
transform 1 0 4704 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_69
timestamp 1698431365
transform 1 0 9072 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_71
timestamp 1698431365
transform 1 0 9296 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_88
timestamp 1698431365
transform 1 0 11200 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_104
timestamp 1698431365
transform 1 0 12992 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_123
timestamp 1698431365
transform 1 0 15120 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_125
timestamp 1698431365
transform 1 0 15344 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_128
timestamp 1698431365
transform 1 0 15680 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_138
timestamp 1698431365
transform 1 0 16800 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_142
timestamp 1698431365
transform 1 0 17248 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_6
timestamp 1698431365
transform 1 0 2016 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_10
timestamp 1698431365
transform 1 0 2464 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_14
timestamp 1698431365
transform 1 0 2912 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_46
timestamp 1698431365
transform 1 0 6496 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_68
timestamp 1698431365
transform 1 0 8960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_76
timestamp 1698431365
transform 1 0 9856 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_120
timestamp 1698431365
transform 1 0 14784 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698431365
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_146
timestamp 1698431365
transform 1 0 17696 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_6
timestamp 1698431365
transform 1 0 2016 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_22
timestamp 1698431365
transform 1 0 3808 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_30
timestamp 1698431365
transform 1 0 4704 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_57
timestamp 1698431365
transform 1 0 7728 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_59
timestamp 1698431365
transform 1 0 7952 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_97
timestamp 1698431365
transform 1 0 12208 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_104
timestamp 1698431365
transform 1 0 12992 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_139
timestamp 1698431365
transform 1 0 16912 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_147
timestamp 1698431365
transform 1 0 17808 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_151
timestamp 1698431365
transform 1 0 18256 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_6
timestamp 1698431365
transform 1 0 2016 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_38
timestamp 1698431365
transform 1 0 5600 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_46
timestamp 1698431365
transform 1 0 6496 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_74
timestamp 1698431365
transform 1 0 9632 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_118
timestamp 1698431365
transform 1 0 14560 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_134
timestamp 1698431365
transform 1 0 16352 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_138
timestamp 1698431365
transform 1 0 16800 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_148
timestamp 1698431365
transform 1 0 17920 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_12
timestamp 1698431365
transform 1 0 2688 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_28
timestamp 1698431365
transform 1 0 4480 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_32
timestamp 1698431365
transform 1 0 4928 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_41
timestamp 1698431365
transform 1 0 5936 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_43
timestamp 1698431365
transform 1 0 6160 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_94
timestamp 1698431365
transform 1 0 11872 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_98
timestamp 1698431365
transform 1 0 12320 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_34
timestamp 1698431365
transform 1 0 5152 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_121
timestamp 1698431365
transform 1 0 14896 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_142
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_102
timestamp 1698431365
transform 1 0 12768 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_112
timestamp 1698431365
transform 1 0 13888 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_144
timestamp 1698431365
transform 1 0 17472 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_6
timestamp 1698431365
transform 1 0 2016 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_22
timestamp 1698431365
transform 1 0 3808 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_30
timestamp 1698431365
transform 1 0 4704 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_34
timestamp 1698431365
transform 1 0 5152 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_74
timestamp 1698431365
transform 1 0 9632 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_82
timestamp 1698431365
transform 1 0 10528 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_103
timestamp 1698431365
transform 1 0 12880 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_135
timestamp 1698431365
transform 1 0 16464 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_139
timestamp 1698431365
transform 1 0 16912 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_150
timestamp 1698431365
transform 1 0 18144 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_8
timestamp 1698431365
transform 1 0 2240 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_12
timestamp 1698431365
transform 1 0 2688 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_28
timestamp 1698431365
transform 1 0 4480 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_32
timestamp 1698431365
transform 1 0 4928 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_37
timestamp 1698431365
transform 1 0 5488 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_94
timestamp 1698431365
transform 1 0 11872 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_102
timestamp 1698431365
transform 1 0 12768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_104
timestamp 1698431365
transform 1 0 12992 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_139
timestamp 1698431365
transform 1 0 16912 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_147
timestamp 1698431365
transform 1 0 17808 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_151
timestamp 1698431365
transform 1 0 18256 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_6
timestamp 1698431365
transform 1 0 2016 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_22
timestamp 1698431365
transform 1 0 3808 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_30
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_34
timestamp 1698431365
transform 1 0 5152 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_36
timestamp 1698431365
transform 1 0 5376 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_11_82
timestamp 1698431365
transform 1 0 10528 0 -1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_114
timestamp 1698431365
transform 1 0 14112 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_130
timestamp 1698431365
transform 1 0 15904 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_150
timestamp 1698431365
transform 1 0 18144 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698431365
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698431365
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_139
timestamp 1698431365
transform 1 0 16912 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_147
timestamp 1698431365
transform 1 0 17808 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_151
timestamp 1698431365
transform 1 0 18256 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_6
timestamp 1698431365
transform 1 0 2016 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698431365
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_6
timestamp 1698431365
transform 1 0 2016 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_22
timestamp 1698431365
transform 1 0 3808 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_30
timestamp 1698431365
transform 1 0 4704 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_89
timestamp 1698431365
transform 1 0 11312 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_139
timestamp 1698431365
transform 1 0 16912 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_14
timestamp 1698431365
transform 1 0 2912 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_18
timestamp 1698431365
transform 1 0 3360 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_23
timestamp 1698431365
transform 1 0 3920 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_31
timestamp 1698431365
transform 1 0 4816 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_35
timestamp 1698431365
transform 1 0 5264 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_41
timestamp 1698431365
transform 1 0 5936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_47
timestamp 1698431365
transform 1 0 6608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_51
timestamp 1698431365
transform 1 0 7056 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_55
timestamp 1698431365
transform 1 0 7504 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_59
timestamp 1698431365
transform 1 0 7952 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_65
timestamp 1698431365
transform 1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_80
timestamp 1698431365
transform 1 0 10304 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_82
timestamp 1698431365
transform 1 0 10528 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_85
timestamp 1698431365
transform 1 0 10864 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_117
timestamp 1698431365
transform 1 0 14448 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_36
timestamp 1698431365
transform 1 0 5376 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_54
timestamp 1698431365
transform 1 0 7392 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_61
timestamp 1698431365
transform 1 0 8176 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_63
timestamp 1698431365
transform 1 0 8400 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_70
timestamp 1698431365
transform 1 0 9184 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_72
timestamp 1698431365
transform 1 0 9408 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_77
timestamp 1698431365
transform 1 0 9968 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_83
timestamp 1698431365
transform 1 0 10640 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_101
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_108
timestamp 1698431365
transform 1 0 13440 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_113
timestamp 1698431365
transform 1 0 14000 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_119
timestamp 1698431365
transform 1 0 14672 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_125
timestamp 1698431365
transform 1 0 15344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_131
timestamp 1698431365
transform 1 0 16016 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_150
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input1
timestamp 1698431365
transform 1 0 7504 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input2
timestamp 1698431365
transform -1 0 18368 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input3
timestamp 1698431365
transform 1 0 2240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input4
timestamp 1698431365
transform -1 0 10864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input5
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input6
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform 1 0 3136 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input8
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform 1 0 4480 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform 1 0 6272 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform 1 0 5488 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input12 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 3808 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 18256 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform 1 0 7616 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 6944 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input16
timestamp 1698431365
transform -1 0 15680 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input17
timestamp 1698431365
transform -1 0 18368 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input18
timestamp 1698431365
transform -1 0 15008 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input19
timestamp 1698431365
transform -1 0 16240 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input20
timestamp 1698431365
transform -1 0 14336 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input21
timestamp 1698431365
transform -1 0 16352 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input22
timestamp 1698431365
transform -1 0 17696 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input23
timestamp 1698431365
transform -1 0 18368 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input24
timestamp 1698431365
transform -1 0 17024 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input25
timestamp 1698431365
transform -1 0 18144 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input26
timestamp 1698431365
transform -1 0 17472 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input27
timestamp 1698431365
transform -1 0 13664 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input28
timestamp 1698431365
transform 1 0 10864 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input29
timestamp 1698431365
transform -1 0 12208 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input30
timestamp 1698431365
transform 1 0 1792 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input31
timestamp 1698431365
transform -1 0 10192 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input32
timestamp 1698431365
transform 1 0 5600 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input33
timestamp 1698431365
transform -1 0 8960 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input34
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input35
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input36
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output37 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 3584 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_3  output38 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 6944 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_4  output39
timestamp 1698431365
transform -1 0 5152 0 1 15680
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_17 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 18592 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_18
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 18592 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_19
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 18592 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_20
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 18592 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_21
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 18592 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_22
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 18592 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_23
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 18592 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_24
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 18592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_25
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 18592 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_26
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 18592 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_27
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 18592 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_28
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 18592 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_29
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 18592 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_30
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 18592 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_31
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 18592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_32
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 18592 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_33
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 18592 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_34 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_35
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_36
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_37
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_38
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_39
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_40
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_41
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_42
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_43
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_44
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_45
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_46
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_47
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_48
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_49
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_50
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_51
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_52
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_53
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_54
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_55
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_56
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_57
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_58
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_59
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_60
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_61
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_62
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_63
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_64
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_65
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_66
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_67
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_68
timestamp 1698431365
transform 1 0 5152 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_69
timestamp 1698431365
transform 1 0 8960 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_70
timestamp 1698431365
transform 1 0 12768 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_71
timestamp 1698431365
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_40 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18144 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_41
timestamp 1698431365
transform -1 0 14000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_42
timestamp 1698431365
transform -1 0 6608 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_43
timestamp 1698431365
transform -1 0 2016 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_44
timestamp 1698431365
transform -1 0 2016 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_45
timestamp 1698431365
transform -1 0 3360 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_46
timestamp 1698431365
transform -1 0 2688 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_47
timestamp 1698431365
transform -1 0 2016 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_48
timestamp 1698431365
transform -1 0 2016 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_49
timestamp 1698431365
transform -1 0 11984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_50
timestamp 1698431365
transform -1 0 10640 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_51
timestamp 1698431365
transform -1 0 13440 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_52
timestamp 1698431365
transform -1 0 17248 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_53
timestamp 1698431365
transform 1 0 17920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_54
timestamp 1698431365
transform 1 0 17472 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_55
timestamp 1698431365
transform -1 0 15344 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_56
timestamp 1698431365
transform -1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_57
timestamp 1698431365
transform -1 0 3920 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_58
timestamp 1698431365
transform -1 0 9968 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_59
timestamp 1698431365
transform -1 0 14672 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_60
timestamp 1698431365
transform -1 0 7392 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_61
timestamp 1698431365
transform 1 0 16128 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_62
timestamp 1698431365
transform -1 0 17696 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_63
timestamp 1698431365
transform -1 0 2016 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_64
timestamp 1698431365
transform -1 0 2016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_65
timestamp 1698431365
transform -1 0 8624 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_66
timestamp 1698431365
transform -1 0 5936 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_67
timestamp 1698431365
transform -1 0 2016 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_68
timestamp 1698431365
transform -1 0 2688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_69
timestamp 1698431365
transform -1 0 16016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  wishbone_register_70
timestamp 1698431365
transform 1 0 8512 0 1 15680
box -86 -86 534 870
<< labels >>
flabel metal2 s 2688 19200 2800 20000 0 FreeSans 448 90 0 0 reg_q_o
port 0 nsew signal tristate
flabel metal4 s 3340 3076 3660 16524 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 7652 3076 7972 16524 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 11964 3076 12284 16524 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 16276 3076 16596 16524 0 FreeSans 1280 90 0 0 vdd
port 1 nsew power bidirectional
flabel metal4 s 5496 3076 5816 16524 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 9808 3076 10128 16524 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 14120 3076 14440 16524 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal4 s 18432 3076 18752 16524 0 FreeSans 1280 90 0 0 vss
port 2 nsew ground bidirectional
flabel metal3 s 0 12096 800 12208 0 FreeSans 448 0 0 0 wb_clk_i
port 3 nsew signal input
flabel metal2 s 7392 19200 7504 20000 0 FreeSans 448 90 0 0 wb_rst_i
port 4 nsew signal input
flabel metal2 s 4704 19200 4816 20000 0 FreeSans 448 90 0 0 wbs_ack_o
port 5 nsew signal tristate
flabel metal2 s 18816 0 18928 800 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 6 nsew signal input
flabel metal2 s 0 0 112 800 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 7 nsew signal input
flabel metal2 s 10080 0 10192 800 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 8 nsew signal input
flabel metal2 s 672 0 784 800 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 9 nsew signal input
flabel metal2 s 1344 0 1456 800 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 10 nsew signal input
flabel metal2 s 3360 0 3472 800 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 11 nsew signal input
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 12 nsew signal input
flabel metal2 s 4704 0 4816 800 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 13 nsew signal input
flabel metal2 s 6720 0 6832 800 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 14 nsew signal input
flabel metal2 s 5376 0 5488 800 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 15 nsew signal input
flabel metal2 s 4032 0 4144 800 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 16 nsew signal input
flabel metal2 s 17472 0 17584 800 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 17 nsew signal input
flabel metal2 s 8064 0 8176 800 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 18 nsew signal input
flabel metal2 s 7392 0 7504 800 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 19 nsew signal input
flabel metal2 s 14112 0 14224 800 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 20 nsew signal input
flabel metal3 s 19200 8736 20000 8848 0 FreeSans 448 0 0 0 wbs_adr_i[23]
port 21 nsew signal input
flabel metal2 s 13440 0 13552 800 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 22 nsew signal input
flabel metal2 s 15456 0 15568 800 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 23 nsew signal input
flabel metal2 s 12768 0 12880 800 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 24 nsew signal input
flabel metal2 s 14784 0 14896 800 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 25 nsew signal input
flabel metal3 s 19200 7392 20000 7504 0 FreeSans 448 0 0 0 wbs_adr_i[28]
port 26 nsew signal input
flabel metal3 s 19200 8064 20000 8176 0 FreeSans 448 0 0 0 wbs_adr_i[29]
port 27 nsew signal input
flabel metal2 s 18144 0 18256 800 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 28 nsew signal input
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 29 nsew signal input
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 30 nsew signal input
flabel metal2 s 12096 0 12208 800 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 31 nsew signal input
flabel metal2 s 10752 0 10864 800 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 32 nsew signal input
flabel metal2 s 11424 0 11536 800 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 33 nsew signal input
flabel metal2 s 2016 0 2128 800 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 34 nsew signal input
flabel metal2 s 9408 0 9520 800 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 35 nsew signal input
flabel metal2 s 6048 0 6160 800 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 36 nsew signal input
flabel metal2 s 8736 0 8848 800 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 37 nsew signal input
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 wbs_cyc_i
port 38 nsew signal input
flabel metal2 s 10752 19200 10864 20000 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 39 nsew signal input
flabel metal3 s 19200 1344 20000 1456 0 FreeSans 448 0 0 0 wbs_dat_i[10]
port 40 nsew signal input
flabel metal3 s 19200 2016 20000 2128 0 FreeSans 448 0 0 0 wbs_dat_i[11]
port 41 nsew signal input
flabel metal3 s 19200 2688 20000 2800 0 FreeSans 448 0 0 0 wbs_dat_i[12]
port 42 nsew signal input
flabel metal3 s 19200 3360 20000 3472 0 FreeSans 448 0 0 0 wbs_dat_i[13]
port 43 nsew signal input
flabel metal3 s 19200 4032 20000 4144 0 FreeSans 448 0 0 0 wbs_dat_i[14]
port 44 nsew signal input
flabel metal3 s 19200 4704 20000 4816 0 FreeSans 448 0 0 0 wbs_dat_i[15]
port 45 nsew signal input
flabel metal3 s 19200 5376 20000 5488 0 FreeSans 448 0 0 0 wbs_dat_i[16]
port 46 nsew signal input
flabel metal3 s 19200 6048 20000 6160 0 FreeSans 448 0 0 0 wbs_dat_i[17]
port 47 nsew signal input
flabel metal3 s 19200 6720 20000 6832 0 FreeSans 448 0 0 0 wbs_dat_i[18]
port 48 nsew signal input
flabel metal3 s 19200 19488 20000 19600 0 FreeSans 448 0 0 0 wbs_dat_i[19]
port 49 nsew signal input
flabel metal3 s 19200 0 20000 112 0 FreeSans 448 0 0 0 wbs_dat_i[1]
port 50 nsew signal input
flabel metal3 s 19200 672 20000 784 0 FreeSans 448 0 0 0 wbs_dat_i[20]
port 51 nsew signal input
flabel metal3 s 19200 10752 20000 10864 0 FreeSans 448 0 0 0 wbs_dat_i[21]
port 52 nsew signal input
flabel metal3 s 19200 10080 20000 10192 0 FreeSans 448 0 0 0 wbs_dat_i[22]
port 53 nsew signal input
flabel metal3 s 19200 9408 20000 9520 0 FreeSans 448 0 0 0 wbs_dat_i[23]
port 54 nsew signal input
flabel metal3 s 19200 11424 20000 11536 0 FreeSans 448 0 0 0 wbs_dat_i[24]
port 55 nsew signal input
flabel metal3 s 19200 13440 20000 13552 0 FreeSans 448 0 0 0 wbs_dat_i[25]
port 56 nsew signal input
flabel metal3 s 19200 12768 20000 12880 0 FreeSans 448 0 0 0 wbs_dat_i[26]
port 57 nsew signal input
flabel metal3 s 19200 12096 20000 12208 0 FreeSans 448 0 0 0 wbs_dat_i[27]
port 58 nsew signal input
flabel metal3 s 19200 14112 20000 14224 0 FreeSans 448 0 0 0 wbs_dat_i[28]
port 59 nsew signal input
flabel metal3 s 19200 16128 20000 16240 0 FreeSans 448 0 0 0 wbs_dat_i[29]
port 60 nsew signal input
flabel metal3 s 19200 15456 20000 15568 0 FreeSans 448 0 0 0 wbs_dat_i[2]
port 61 nsew signal input
flabel metal3 s 19200 14784 20000 14896 0 FreeSans 448 0 0 0 wbs_dat_i[30]
port 62 nsew signal input
flabel metal3 s 19200 16800 20000 16912 0 FreeSans 448 0 0 0 wbs_dat_i[31]
port 63 nsew signal input
flabel metal3 s 19200 18816 20000 18928 0 FreeSans 448 0 0 0 wbs_dat_i[3]
port 64 nsew signal input
flabel metal3 s 19200 18144 20000 18256 0 FreeSans 448 0 0 0 wbs_dat_i[4]
port 65 nsew signal input
flabel metal3 s 19200 17472 20000 17584 0 FreeSans 448 0 0 0 wbs_dat_i[5]
port 66 nsew signal input
flabel metal2 s 672 19200 784 20000 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 67 nsew signal input
flabel metal2 s 1344 19200 1456 20000 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 68 nsew signal input
flabel metal2 s 0 19200 112 20000 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 69 nsew signal input
flabel metal2 s 2016 19200 2128 20000 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 70 nsew signal input
flabel metal2 s 4032 19200 4144 20000 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 71 nsew signal tristate
flabel metal2 s 11424 19200 11536 20000 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 72 nsew signal tristate
flabel metal2 s 10080 19200 10192 20000 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 73 nsew signal tristate
flabel metal2 s 12768 19200 12880 20000 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 74 nsew signal tristate
flabel metal2 s 16128 19200 16240 20000 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 75 nsew signal tristate
flabel metal2 s 18816 19200 18928 20000 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 76 nsew signal tristate
flabel metal2 s 18144 19200 18256 20000 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 77 nsew signal tristate
flabel metal2 s 14784 19200 14896 20000 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 78 nsew signal tristate
flabel metal2 s 12096 19200 12208 20000 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 79 nsew signal tristate
flabel metal2 s 3360 19200 3472 20000 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 80 nsew signal tristate
flabel metal2 s 9408 19200 9520 20000 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 81 nsew signal tristate
flabel metal2 s 17472 19200 17584 20000 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 82 nsew signal tristate
flabel metal2 s 14112 19200 14224 20000 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 83 nsew signal tristate
flabel metal2 s 6720 19200 6832 20000 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 84 nsew signal tristate
flabel metal2 s 19488 19200 19600 20000 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 85 nsew signal tristate
flabel metal2 s 16800 19200 16912 20000 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 86 nsew signal tristate
flabel metal3 s 0 14112 800 14224 0 FreeSans 448 0 0 0 wbs_dat_o[24]
port 87 nsew signal tristate
flabel metal3 s 0 15456 800 15568 0 FreeSans 448 0 0 0 wbs_dat_o[25]
port 88 nsew signal tristate
flabel metal2 s 8064 19200 8176 20000 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 89 nsew signal tristate
flabel metal2 s 5376 19200 5488 20000 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 90 nsew signal tristate
flabel metal3 s 0 5376 800 5488 0 FreeSans 448 0 0 0 wbs_dat_o[28]
port 91 nsew signal tristate
flabel metal3 s 0 4704 800 4816 0 FreeSans 448 0 0 0 wbs_dat_o[29]
port 92 nsew signal tristate
flabel metal2 s 13440 19200 13552 20000 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 93 nsew signal tristate
flabel metal2 s 15456 19200 15568 20000 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 94 nsew signal tristate
flabel metal2 s 8736 19200 8848 20000 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 95 nsew signal tristate
flabel metal2 s 6048 19200 6160 20000 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 96 nsew signal tristate
flabel metal3 s 0 14784 800 14896 0 FreeSans 448 0 0 0 wbs_dat_o[4]
port 97 nsew signal tristate
flabel metal3 s 0 11424 800 11536 0 FreeSans 448 0 0 0 wbs_dat_o[5]
port 98 nsew signal tristate
flabel metal3 s 0 4032 800 4144 0 FreeSans 448 0 0 0 wbs_dat_o[6]
port 99 nsew signal tristate
flabel metal3 s 0 7392 800 7504 0 FreeSans 448 0 0 0 wbs_dat_o[7]
port 100 nsew signal tristate
flabel metal3 s 0 10080 800 10192 0 FreeSans 448 0 0 0 wbs_dat_o[8]
port 101 nsew signal tristate
flabel metal3 s 0 13440 800 13552 0 FreeSans 448 0 0 0 wbs_dat_o[9]
port 102 nsew signal tristate
flabel metal3 s 0 19488 800 19600 0 FreeSans 448 0 0 0 wbs_sel_i[0]
port 103 nsew signal input
flabel metal3 s 0 18816 800 18928 0 FreeSans 448 0 0 0 wbs_sel_i[1]
port 104 nsew signal input
flabel metal3 s 0 18144 800 18256 0 FreeSans 448 0 0 0 wbs_sel_i[2]
port 105 nsew signal input
flabel metal3 s 0 17472 800 17584 0 FreeSans 448 0 0 0 wbs_sel_i[3]
port 106 nsew signal input
flabel metal3 s 0 8064 800 8176 0 FreeSans 448 0 0 0 wbs_stb_i
port 107 nsew signal input
flabel metal3 s 0 10752 800 10864 0 FreeSans 448 0 0 0 wbs_we_i
port 108 nsew signal input
rlabel metal1 9968 16464 9968 16464 0 vdd
rlabel via1 10048 15680 10048 15680 0 vss
rlabel metal2 8344 9856 8344 9856 0 _00_
rlabel metal2 8344 11368 8344 11368 0 _01_
rlabel metal2 6104 9296 6104 9296 0 _02_
rlabel metal2 6104 11648 6104 11648 0 _03_
rlabel metal3 11312 6664 11312 6664 0 _04_
rlabel metal2 12936 6720 12936 6720 0 _05_
rlabel metal2 12712 8736 12712 8736 0 _06_
rlabel metal2 13384 8960 13384 8960 0 _07_
rlabel metal2 14448 7448 14448 7448 0 _08_
rlabel metal2 10360 6552 10360 6552 0 _09_
rlabel metal2 9912 10080 9912 10080 0 _10_
rlabel metal3 10304 10360 10304 10360 0 _11_
rlabel metal3 9016 5096 9016 5096 0 _12_
rlabel metal2 10360 5432 10360 5432 0 _13_
rlabel metal2 9688 5712 9688 5712 0 _14_
rlabel metal2 11032 6440 11032 6440 0 _15_
rlabel metal2 11144 6440 11144 6440 0 _16_
rlabel metal2 13776 9688 13776 9688 0 _17_
rlabel metal2 13440 9800 13440 9800 0 _18_
rlabel metal2 7616 9800 7616 9800 0 _19_
rlabel metal2 12488 10248 12488 10248 0 _20_
rlabel metal2 10360 9688 10360 9688 0 _21_
rlabel metal2 9688 9632 9688 9632 0 _22_
rlabel metal2 10472 9744 10472 9744 0 clknet_0_wb_clk_i
rlabel metal2 5656 8680 5656 8680 0 clknet_1_0__leaf_wb_clk_i
rlabel metal2 6216 13272 6216 13272 0 clknet_1_1__leaf_wb_clk_i
rlabel metal2 8008 15484 8008 15484 0 net1
rlabel metal3 7504 6664 7504 6664 0 net10
rlabel metal2 5992 4704 5992 4704 0 net11
rlabel metal3 4312 4032 4312 4032 0 net12
rlabel metal2 10248 5208 10248 5208 0 net13
rlabel metal2 8120 3332 8120 3332 0 net14
rlabel metal2 7504 5096 7504 5096 0 net15
rlabel metal2 15176 4648 15176 4648 0 net16
rlabel metal2 17976 7196 17976 7196 0 net17
rlabel metal2 14504 4704 14504 4704 0 net18
rlabel metal2 14616 5208 14616 5208 0 net19
rlabel metal2 17864 5320 17864 5320 0 net2
rlabel metal2 13608 5768 13608 5768 0 net20
rlabel metal2 15848 3752 15848 3752 0 net21
rlabel metal2 17192 8176 17192 8176 0 net22
rlabel metal2 14728 8568 14728 8568 0 net23
rlabel metal2 16520 4760 16520 4760 0 net24
rlabel metal2 17640 3808 17640 3808 0 net25
rlabel metal2 16968 3584 16968 3584 0 net26
rlabel metal2 12824 7728 12824 7728 0 net27
rlabel metal2 11368 6272 11368 6272 0 net28
rlabel metal2 11704 6216 11704 6216 0 net29
rlabel metal2 2856 5992 2856 5992 0 net3
rlabel metal2 2296 3920 2296 3920 0 net30
rlabel metal2 8848 5992 8848 5992 0 net31
rlabel metal3 6608 5992 6608 5992 0 net32
rlabel metal2 7784 5768 7784 5768 0 net33
rlabel metal2 11592 11704 11592 11704 0 net34
rlabel metal2 12712 7280 12712 7280 0 net35
rlabel metal2 2072 10472 2072 10472 0 net36
rlabel metal2 3192 13048 3192 13048 0 net37
rlabel metal3 7896 16072 7896 16072 0 net38
rlabel metal2 9016 12768 9016 12768 0 net39
rlabel metal2 10360 3332 10360 3332 0 net4
rlabel metal2 17696 15960 17696 15960 0 net40
rlabel metal2 13608 15960 13608 15960 0 net41
rlabel metal2 6216 15512 6216 15512 0 net42
rlabel metal3 1246 14840 1246 14840 0 net43
rlabel metal3 1246 11480 1246 11480 0 net44
rlabel metal3 1918 4088 1918 4088 0 net45
rlabel metal3 1582 7448 1582 7448 0 net46
rlabel metal3 1246 10136 1246 10136 0 net47
rlabel metal3 1246 13496 1246 13496 0 net48
rlabel metal2 11592 15960 11592 15960 0 net49
rlabel metal2 2072 5712 2072 5712 0 net5
rlabel metal2 10248 15960 10248 15960 0 net50
rlabel metal2 13160 16744 13160 16744 0 net51
rlabel metal3 16576 15960 16576 15960 0 net52
rlabel metal2 18200 16128 18200 16128 0 net53
rlabel metal2 17752 15624 17752 15624 0 net54
rlabel metal2 14952 15960 14952 15960 0 net55
rlabel metal2 12376 16744 12376 16744 0 net56
rlabel metal2 3696 15512 3696 15512 0 net57
rlabel metal2 9576 15960 9576 15960 0 net58
rlabel metal2 14280 15960 14280 15960 0 net59
rlabel metal2 7336 5992 7336 5992 0 net6
rlabel metal2 7112 16800 7112 16800 0 net60
rlabel metal3 17976 15848 17976 15848 0 net61
rlabel metal2 17416 16352 17416 16352 0 net62
rlabel metal3 1246 14168 1246 14168 0 net63
rlabel metal3 1246 15512 1246 15512 0 net64
rlabel metal2 8232 15512 8232 15512 0 net65
rlabel metal2 5544 15512 5544 15512 0 net66
rlabel metal3 1246 5432 1246 5432 0 net67
rlabel metal3 1582 4760 1582 4760 0 net68
rlabel metal2 15624 15960 15624 15960 0 net69
rlabel metal3 7168 3416 7168 3416 0 net7
rlabel metal2 8792 17626 8792 17626 0 net70
rlabel metal2 5880 11928 5880 11928 0 net71
rlabel metal2 2968 4928 2968 4928 0 net8
rlabel metal2 4984 4200 4984 4200 0 net9
rlabel metal2 2744 17738 2744 17738 0 reg_q_o
rlabel metal3 5824 11368 5824 11368 0 wb_clk_i
rlabel metal2 7560 16072 7560 16072 0 wb_rst_i
rlabel metal3 5376 16296 5376 16296 0 wbs_ack_o
rlabel metal2 18200 4368 18200 4368 0 wbs_adr_i[0]
rlabel metal2 2408 3864 2408 3864 0 wbs_adr_i[10]
rlabel metal2 10192 2856 10192 2856 0 wbs_adr_i[11]
rlabel metal2 1736 5040 1736 5040 0 wbs_adr_i[12]
rlabel metal2 1736 3976 1736 3976 0 wbs_adr_i[13]
rlabel metal2 3584 3640 3584 3640 0 wbs_adr_i[14]
rlabel metal2 2744 2142 2744 2142 0 wbs_adr_i[15]
rlabel metal2 4816 4200 4816 4200 0 wbs_adr_i[16]
rlabel metal2 6720 3080 6720 3080 0 wbs_adr_i[17]
rlabel metal2 5656 4256 5656 4256 0 wbs_adr_i[18]
rlabel metal2 4256 4200 4256 4200 0 wbs_adr_i[19]
rlabel metal2 17920 4312 17920 4312 0 wbs_adr_i[1]
rlabel metal2 8120 854 8120 854 0 wbs_adr_i[20]
rlabel metal2 7504 2520 7504 2520 0 wbs_adr_i[21]
rlabel metal2 14168 1302 14168 1302 0 wbs_adr_i[22]
rlabel metal2 18200 8904 18200 8904 0 wbs_adr_i[23]
rlabel metal2 13776 2296 13776 2296 0 wbs_adr_i[24]
rlabel metal2 15568 4200 15568 4200 0 wbs_adr_i[25]
rlabel metal3 13496 3416 13496 3416 0 wbs_adr_i[26]
rlabel metal2 16072 3472 16072 3472 0 wbs_adr_i[27]
rlabel metal3 18522 7448 18522 7448 0 wbs_adr_i[28]
rlabel metal3 18746 8120 18746 8120 0 wbs_adr_i[29]
rlabel metal3 17472 4312 17472 4312 0 wbs_adr_i[2]
rlabel metal2 17976 3192 17976 3192 0 wbs_adr_i[30]
rlabel metal2 17192 3472 17192 3472 0 wbs_adr_i[31]
rlabel metal2 12152 2058 12152 2058 0 wbs_adr_i[3]
rlabel metal2 10920 3528 10920 3528 0 wbs_adr_i[4]
rlabel metal3 11704 3528 11704 3528 0 wbs_adr_i[5]
rlabel metal2 1960 4312 1960 4312 0 wbs_adr_i[6]
rlabel metal2 9912 3416 9912 3416 0 wbs_adr_i[7]
rlabel metal2 5992 2296 5992 2296 0 wbs_adr_i[8]
rlabel metal2 8792 2058 8792 2058 0 wbs_adr_i[9]
rlabel metal2 10920 16072 10920 16072 0 wbs_dat_i[0]
rlabel metal2 4088 17738 4088 17738 0 wbs_dat_o[0]
rlabel metal3 1246 8120 1246 8120 0 wbs_stb_i
rlabel metal2 1848 11088 1848 11088 0 wbs_we_i
<< properties >>
string FIXED_BBOX 0 0 20000 20000
<< end >>
